library ieee;
library work;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use work.arrayAsAliasTrimmers.all;
use work.types.all;
use work.runtime.all;
use work.IOShuvalkin.all;
use work.bincompl.all;
library unisim;
library UNISIM;
entity proc_TopMain is
port (clk : in std_logic;
      rst : in std_logic
      ;
      
      -- input signals
      reset_ena     : in std_logic; 
       
      outp_rdy_ena     : in std_logic; 
       
      outpVars_rdy_ena     : in std_logic; 
       
      outp1_rdy_ena     : in std_logic; 
       
      inp_data     : in recinp2; 
       
      inp_ena     : in std_logic
      ;
      
      -- -- output signals
      reset_rdy_ena     : out std_logic; 
       
      outpVars_data     : out recoutpVars; 
       
      outpVars_ena     : out std_logic; 
       
      outp1_data     : out recoutp; 
       
      outp1_ena     : out std_logic; 
       
      outp_data     : out recoutp; 
       
      outp_ena     : out std_logic; 
       
      inp_rdy_ena     : out std_logic);
end entity;
architecture rtl of proc_TopMain is 
signal cycleNum : integer;
signal defihscl0000035 : std_logic_vector (0 downto 0) := std_logic_vector'(B"1");
signal endofoutphscl0000036 : std_logic_vector (0 downto 0) :=  conv_std_logic_vector
                                                               (0,  1);
signal endofoutp1hscl0000037 : std_logic_vector (0 downto 0) :=  conv_std_logic_vector
                                                                (0,  1);
signal h0_elseTransactionhscl0000038 : std_logic_vector (0 downto 0) := (0 => '0');
signal h1_elseTransactionhscl0000039 : std_logic_vector (0 downto 0) := (0 => '0');
signal h1_then_l_elseTransactionhscl000003a : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h1_then_l_then_lastHappened0hscl000003b : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h1_then_l_then_lastHappened1hscl000003c : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h1_then_l_then_lastHappened2hscl000003d : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h1_then_l_then_p2_elseTransactionhscl000003e : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h1_then_leftHappenedhscl000003f : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h2_elseTransactionhscl000003g : std_logic_vector (0 downto 0) := (0 => '0');
signal h2_else_elseTransactionhscl000003h : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h3_elseTransactionhscl000003i : std_logic_vector (0 downto 0) := (0 => '0');
signal h3_else_elseTransactionhscl000003j : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h4_elseTransactionhscl000003k : std_logic_vector (0 downto 0) := (0 => '0');
signal h5_elseTransactionhscl000003l : std_logic_vector (0 downto 0) := (0 => '0');
signal h5_then_elseTransactionhscl000003m : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h5_then_then_elseTransactionhscl000003n : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h5_then_then_else_l_lastHappened0hscl000003o : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h5_then_then_else_l_lastHappened1hscl000003p : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h5_then_then_else_l_lastHappened2hscl000003q : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h5_then_then_else_l_p0_elseTransactionhscl000003r : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h5_then_then_else_leftHappenedhscl000003s : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h5_then_then_then_l_lastHappened0hscl000003t : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h5_then_then_then_l_lastHappened1hscl000003u : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h5_then_then_then_l_lastHappened2hscl000003v : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h5_then_then_then_leftHappenedhscl000003w : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h6_elseTransactionhscl000003x : std_logic_vector (0 downto 0) := (0 => '0');
signal h7_elseTransactionhscl000003y : std_logic_vector (0 downto 0) := (0 => '0');
signal h7_then_lastHappened0hscl000003z : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_lastHappened1hscl0000040 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p0_elseTransactionhscl0000041 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p0_then_lastHappened0hscl0000042 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p0_then_lastHappened1hscl0000043 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p0_then_lastHappened2hscl0000044 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p0_then_p2_lastHappened0hscl0000045 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p0_then_p2_lastHappened1hscl0000046 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p0_then_p2_lastHappened2hscl0000047 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p0_then_p2_p2_elseTransactionhscl0000048 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_elseTransactionhscl0000049 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened0hscl000004a : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened1hscl000004b : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened10hscl000004c : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened11hscl000004d : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened12hscl000004e : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened13hscl000004f : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened14hscl000004g : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened15hscl000004h : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened16hscl000004i : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened17hscl000004j : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened18hscl000004k : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened19hscl000004l : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened2hscl000004m : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened20hscl000004n : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened21hscl000004o : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened22hscl000004p : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened23hscl000004q : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened24hscl000004r : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened25hscl000004s : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened26hscl000004t : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened27hscl000004u : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened28hscl000004v : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened29hscl000004w : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened3hscl000004x : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened30hscl000004y : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened31hscl000004z : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened32hscl0000050 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened33hscl0000051 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened34hscl0000052 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened35hscl0000053 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened36hscl0000054 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened37hscl0000055 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened38hscl0000056 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened39hscl0000057 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened4hscl0000058 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened40hscl0000059 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened41hscl000005a : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened42hscl000005b : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened43hscl000005c : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened44hscl000005d : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened45hscl000005e : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened46hscl000005f : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened47hscl000005g : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened48hscl000005h : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened49hscl000005i : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened5hscl000005j : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened50hscl000005k : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened51hscl000005l : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened52hscl000005m : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened53hscl000005n : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened54hscl000005o : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened55hscl000005p : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened56hscl000005q : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened57hscl000005r : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened58hscl000005s : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened59hscl000005t : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened6hscl000005u : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened60hscl000005v : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened61hscl000005w : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened62hscl000005x : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened63hscl000005y : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened64hscl000005z : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened7hscl0000060 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened8hscl0000061 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal h7_then_p1_then_lastHappened9hscl0000062 : std_logic_vector (0 downto 0)
 := (0 => '0');
signal ihscl0000063 :  std_logic_vector (10-1 downto 0) :=  conv_std_logic_vector
                                                           (0,  10);
signal icoefmulthscl0000064 : arrticoefmult1(0 to 63);
signal sumshscl0000065 : arrtsums1(0 to 63);
signal sumsqshscl0000066 : arrtsumsqs1(0 to 63);
signal varLefthscl0000067 : arrtvarLeft1(0 to 63);
signal varLeft1hscl0000068 : arrtvarLeft11(0 to 63);
signal varLeft2hscl0000069 : arrtvarLeft11(0 to 63);
signal varRighthscl000006a : arrtvarLeft1(0 to 63);
signal varRight1hscl000006b : arrtvarRight11(0 to 63);
signal varRight2hscl000006c : arrtvarRight11(0 to 63);
signal handlerForVar_rdyhscl000001g_ena : std_logic;
signal handlerForVarRCut_rdyhscl000001e_ena : std_logic;
signal handlerForVarRCuthscl000001h_data : recinp;
signal handlerForVarRCuthscl000001h_ena : std_logic;
signal handlerForVarhscl000001f_data : recinp;
signal handlerForVarhscl000001f_ena : std_logic;
signal h7_then_p1_then_enablehscl0000034_ena : std_logic;
signal h7_then_p1_thenEnablehscl0000033_ena : std_logic;
signal h7_then_p1_elseEnablehscl0000032_ena : std_logic;
signal h7_then_p0_then_p2_p2_thenEnablehscl0000031_ena : std_logic;
signal h7_then_p0_then_p2_p2_elseEnablehscl0000030_ena : std_logic;
signal h7_then_p0_then_p2_enablehscl000002z_ena : std_logic;
signal h7_then_p0_then_enablehscl000002y_ena : std_logic;
signal h7_then_p0_thenEnablehscl000002x_ena : std_logic;
signal h7_then_p0_elseEnablehscl000002w_ena : std_logic;
signal h7_then_enablehscl000002v_ena : std_logic;
signal h7_thenEnablehscl000002u_ena : std_logic;
signal h7_elseEnablehscl000002t_ena : std_logic;
signal h6_thenEnablehscl000002s_ena : std_logic;
signal h6_elseEnablehscl000002r_ena : std_logic;
signal h5_then_then_then_rightEnablehscl000002q_ena : std_logic;
signal h5_then_then_then_l_enablehscl000002p_ena : std_logic;
signal h5_then_then_then_enablehscl000002o_ena : std_logic;
signal h5_then_then_thenEnablehscl000002n_ena : std_logic;
signal h5_then_then_else_rightEnablehscl000002m_ena : std_logic;
signal h5_then_then_else_l_p0_thenEnablehscl000002l_ena : std_logic;
signal h5_then_then_else_l_p0_elseEnablehscl000002k_ena : std_logic;
signal h5_then_then_else_l_enablehscl000002j_ena : std_logic;
signal h5_then_then_else_enablehscl000002i_ena : std_logic;
signal h5_then_then_elseEnablehscl000002h_ena : std_logic;
signal h5_then_thenEnablehscl000002g_ena : std_logic;
signal h5_then_elseEnablehscl000002f_ena : std_logic;
signal h5_thenEnablehscl000002e_ena : std_logic;
signal h5_elseEnablehscl000002d_ena : std_logic;
signal h4_thenEnablehscl000002c_ena : std_logic;
signal h4_elseEnablehscl000002b_ena : std_logic;
signal h3_thenEnablehscl000002a_ena : std_logic;
signal h3_else_thenEnablehscl0000029_ena : std_logic;
signal h3_else_elseEnablehscl0000028_ena : std_logic;
signal h3_elseEnablehscl0000027_ena : std_logic;
signal h2_thenEnablehscl0000026_ena : std_logic;
signal h2_else_thenEnablehscl0000025_ena : std_logic;
signal h2_else_elseEnablehscl0000024_ena : std_logic;
signal h2_elseEnablehscl0000023_ena : std_logic;
signal h1s_finish4_rdyhscl0000022_ena : std_logic;
signal h1s_finish4hscl0000021_ena : std_logic;
signal h1sT_finish_rdyhscl0000020_ena : std_logic;
signal h1sT_finish4_rdyhscl000001z_ena : std_logic;
signal h1sT_finish4hscl000001y_data : recinp2;
signal h1sT_finish4hscl000001y_ena : std_logic;
signal h1sT_finishhscl000001x_data : recinp2;
signal h1sT_finishhscl000001x_ena : std_logic;
signal h1sTT_finish_rdyhscl000001w_ena : std_logic;
signal h1sTT_finish4_rdyhscl000001v_ena : std_logic;
signal h1sTT_finish4hscl000001u_data : recinp2;
signal h1sTT_finish4hscl000001u_ena : std_logic;
signal h1sTT_finishhscl000001t_data : recinp2;
signal h1sTT_finishhscl000001t_ena : std_logic;
signal h1sTTE_finish_rdyhscl0000014_ena : std_logic;
signal h1sTTE_finish4_rdyhscl000001a_ena : std_logic;
signal h1sTTE_finish4hscl000001d_data : recinp2;
signal h1sTTE_finish4hscl000001d_ena : std_logic;
signal h1sTTE_finish3_rdyhscl000001c_ena : std_logic;
signal h1sTTE_finish3hscl000001b_data : recinp2;
signal h1sTTE_finish3hscl000001b_ena : std_logic;
signal h1sTTE_finish2_rdyhscl0000017_ena : std_logic;
signal h1sTTE_finish2hscl0000019_data : recinp2;
signal h1sTTE_finish2hscl0000019_ena : std_logic;
signal h1sTTE_finish1_rdyhscl0000012_ena : std_logic;
signal h1sTTE_finish1hscl0000015_data : recinp2;
signal h1sTTE_finish1hscl0000015_ena : std_logic;
signal h1sTTE_finishhscl0000013_data : recinp2;
signal h1sTTE_finishhscl0000013_ena : std_logic;
signal h1_then_rightEnablehscl000001s_ena : std_logic;
signal h1_then_l_then_p2_thenEnablehscl000001r_ena : std_logic;
signal h1_then_l_then_p2_elseEnablehscl000001q_ena : std_logic;
signal h1_then_l_then_enablehscl000001p_ena : std_logic;
signal h1_then_l_thenEnablehscl000001o_ena : std_logic;
signal h1_then_l_elseEnablehscl000001n_ena : std_logic;
signal h1_then_enablehscl000001m_ena : std_logic;
signal h1_thenEnablehscl000001l_ena : std_logic;
signal h1_elseEnablehscl000001k_ena : std_logic;
signal h0_thenEnablehscl000001j_ena : std_logic;
signal h0_elseEnablehscl000001i_ena : std_logic;
signal Pipe_h1sTTE0BufFull_rdyhscl0000016_ena : std_logic;
signal Pipe_h1sTTE0BufFullhscl0000018_ena : std_logic;
file defitrace : char_file open write_mode is "Top.Maindefi.trace";
file endofoutptrace : char_file open write_mode is "Top.Mainendofoutp.trace";
file endofoutp1trace : char_file open write_mode is "Top.Mainendofoutp1.trace";
file h0_elseTransactiontrace : char_file open write_mode is "Top.Mainh0_elseTransaction.trace";
file h1_elseTransactiontrace : char_file open write_mode is "Top.Mainh1_elseTransaction.trace";
file h1_then_l_elseTransactiontrace : char_file open write_mode is "Top.Mainh1_then_l_elseTransaction.trace";
file h1_then_l_then_lastHappened0trace : char_file open write_mode is "Top.Mainh1_then_l_then_lastHappened0.trace";
file h1_then_l_then_lastHappened1trace : char_file open write_mode is "Top.Mainh1_then_l_then_lastHappened1.trace";
file h1_then_l_then_lastHappened2trace : char_file open write_mode is "Top.Mainh1_then_l_then_lastHappened2.trace";
file h1_then_l_then_p2_elseTransactiontrace : char_file open write_mode is "Top.Mainh1_then_l_then_p2_elseTransaction.trace";
file h1_then_leftHappenedtrace : char_file open write_mode is "Top.Mainh1_then_leftHappened.trace";
file h2_elseTransactiontrace : char_file open write_mode is "Top.Mainh2_elseTransaction.trace";
file h2_else_elseTransactiontrace : char_file open write_mode is "Top.Mainh2_else_elseTransaction.trace";
file h3_elseTransactiontrace : char_file open write_mode is "Top.Mainh3_elseTransaction.trace";
file h3_else_elseTransactiontrace : char_file open write_mode is "Top.Mainh3_else_elseTransaction.trace";
file h4_elseTransactiontrace : char_file open write_mode is "Top.Mainh4_elseTransaction.trace";
file h5_elseTransactiontrace : char_file open write_mode is "Top.Mainh5_elseTransaction.trace";
file h5_then_elseTransactiontrace : char_file open write_mode is "Top.Mainh5_then_elseTransaction.trace";
file h5_then_then_elseTransactiontrace : char_file open write_mode is "Top.Mainh5_then_then_elseTransaction.trace";
file h5_then_then_else_l_lastHappened0trace : char_file open write_mode is "Top.Mainh5_then_then_else_l_lastHappened0.trace";
file h5_then_then_else_l_lastHappened1trace : char_file open write_mode is "Top.Mainh5_then_then_else_l_lastHappened1.trace";
file h5_then_then_else_l_lastHappened2trace : char_file open write_mode is "Top.Mainh5_then_then_else_l_lastHappened2.trace";
file h5_then_then_else_l_p0_elseTransactiontrace : char_file open write_mode is "Top.Mainh5_then_then_else_l_p0_elseTransaction.trace";
file h5_then_then_else_leftHappenedtrace : char_file open write_mode is "Top.Mainh5_then_then_else_leftHappened.trace";
file h5_then_then_then_l_lastHappened0trace : char_file open write_mode is "Top.Mainh5_then_then_then_l_lastHappened0.trace";
file h5_then_then_then_l_lastHappened1trace : char_file open write_mode is "Top.Mainh5_then_then_then_l_lastHappened1.trace";
file h5_then_then_then_l_lastHappened2trace : char_file open write_mode is "Top.Mainh5_then_then_then_l_lastHappened2.trace";
file h5_then_then_then_leftHappenedtrace : char_file open write_mode is "Top.Mainh5_then_then_then_leftHappened.trace";
file h6_elseTransactiontrace : char_file open write_mode is "Top.Mainh6_elseTransaction.trace";
file h7_elseTransactiontrace : char_file open write_mode is "Top.Mainh7_elseTransaction.trace";
file h7_then_lastHappened0trace : char_file open write_mode is "Top.Mainh7_then_lastHappened0.trace";
file h7_then_lastHappened1trace : char_file open write_mode is "Top.Mainh7_then_lastHappened1.trace";
file h7_then_p0_elseTransactiontrace : char_file open write_mode is "Top.Mainh7_then_p0_elseTransaction.trace";
file h7_then_p0_then_lastHappened0trace : char_file open write_mode is "Top.Mainh7_then_p0_then_lastHappened0.trace";
file h7_then_p0_then_lastHappened1trace : char_file open write_mode is "Top.Mainh7_then_p0_then_lastHappened1.trace";
file h7_then_p0_then_lastHappened2trace : char_file open write_mode is "Top.Mainh7_then_p0_then_lastHappened2.trace";
file h7_then_p0_then_p2_lastHappened0trace : char_file open write_mode is "Top.Mainh7_then_p0_then_p2_lastHappened0.trace";
file h7_then_p0_then_p2_lastHappened1trace : char_file open write_mode is "Top.Mainh7_then_p0_then_p2_lastHappened1.trace";
file h7_then_p0_then_p2_lastHappened2trace : char_file open write_mode is "Top.Mainh7_then_p0_then_p2_lastHappened2.trace";
file h7_then_p0_then_p2_p2_elseTransactiontrace : char_file open write_mode is "Top.Mainh7_then_p0_then_p2_p2_elseTransaction.trace";
file h7_then_p1_elseTransactiontrace : char_file open write_mode is "Top.Mainh7_then_p1_elseTransaction.trace";
file h7_then_p1_then_lastHappened0trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened0.trace";
file h7_then_p1_then_lastHappened1trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened1.trace";
file h7_then_p1_then_lastHappened10trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened10.trace";
file h7_then_p1_then_lastHappened11trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened11.trace";
file h7_then_p1_then_lastHappened12trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened12.trace";
file h7_then_p1_then_lastHappened13trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened13.trace";
file h7_then_p1_then_lastHappened14trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened14.trace";
file h7_then_p1_then_lastHappened15trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened15.trace";
file h7_then_p1_then_lastHappened16trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened16.trace";
file h7_then_p1_then_lastHappened17trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened17.trace";
file h7_then_p1_then_lastHappened18trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened18.trace";
file h7_then_p1_then_lastHappened19trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened19.trace";
file h7_then_p1_then_lastHappened2trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened2.trace";
file h7_then_p1_then_lastHappened20trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened20.trace";
file h7_then_p1_then_lastHappened21trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened21.trace";
file h7_then_p1_then_lastHappened22trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened22.trace";
file h7_then_p1_then_lastHappened23trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened23.trace";
file h7_then_p1_then_lastHappened24trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened24.trace";
file h7_then_p1_then_lastHappened25trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened25.trace";
file h7_then_p1_then_lastHappened26trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened26.trace";
file h7_then_p1_then_lastHappened27trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened27.trace";
file h7_then_p1_then_lastHappened28trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened28.trace";
file h7_then_p1_then_lastHappened29trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened29.trace";
file h7_then_p1_then_lastHappened3trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened3.trace";
file h7_then_p1_then_lastHappened30trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened30.trace";
file h7_then_p1_then_lastHappened31trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened31.trace";
file h7_then_p1_then_lastHappened32trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened32.trace";
file h7_then_p1_then_lastHappened33trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened33.trace";
file h7_then_p1_then_lastHappened34trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened34.trace";
file h7_then_p1_then_lastHappened35trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened35.trace";
file h7_then_p1_then_lastHappened36trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened36.trace";
file h7_then_p1_then_lastHappened37trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened37.trace";
file h7_then_p1_then_lastHappened38trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened38.trace";
file h7_then_p1_then_lastHappened39trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened39.trace";
file h7_then_p1_then_lastHappened4trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened4.trace";
file h7_then_p1_then_lastHappened40trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened40.trace";
file h7_then_p1_then_lastHappened41trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened41.trace";
file h7_then_p1_then_lastHappened42trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened42.trace";
file h7_then_p1_then_lastHappened43trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened43.trace";
file h7_then_p1_then_lastHappened44trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened44.trace";
file h7_then_p1_then_lastHappened45trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened45.trace";
file h7_then_p1_then_lastHappened46trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened46.trace";
file h7_then_p1_then_lastHappened47trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened47.trace";
file h7_then_p1_then_lastHappened48trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened48.trace";
file h7_then_p1_then_lastHappened49trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened49.trace";
file h7_then_p1_then_lastHappened5trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened5.trace";
file h7_then_p1_then_lastHappened50trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened50.trace";
file h7_then_p1_then_lastHappened51trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened51.trace";
file h7_then_p1_then_lastHappened52trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened52.trace";
file h7_then_p1_then_lastHappened53trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened53.trace";
file h7_then_p1_then_lastHappened54trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened54.trace";
file h7_then_p1_then_lastHappened55trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened55.trace";
file h7_then_p1_then_lastHappened56trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened56.trace";
file h7_then_p1_then_lastHappened57trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened57.trace";
file h7_then_p1_then_lastHappened58trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened58.trace";
file h7_then_p1_then_lastHappened59trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened59.trace";
file h7_then_p1_then_lastHappened6trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened6.trace";
file h7_then_p1_then_lastHappened60trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened60.trace";
file h7_then_p1_then_lastHappened61trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened61.trace";
file h7_then_p1_then_lastHappened62trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened62.trace";
file h7_then_p1_then_lastHappened63trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened63.trace";
file h7_then_p1_then_lastHappened64trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened64.trace";
file h7_then_p1_then_lastHappened7trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened7.trace";
file h7_then_p1_then_lastHappened8trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened8.trace";
file h7_then_p1_then_lastHappened9trace : char_file open write_mode is "Top.Mainh7_then_p1_then_lastHappened9.trace";
file itrace : char_file open write_mode is "Top.Maini.trace";
file icoefmulttrace : char_file open write_mode is "Top.Mainicoefmult.trace";
file sumstrace : char_file open write_mode is "Top.Mainsums.trace";
file sumsqstrace : char_file open write_mode is "Top.Mainsumsqs.trace";
file varLefttrace : char_file open write_mode is "Top.MainvarLeft.trace";
file varLeft1trace : char_file open write_mode is "Top.MainvarLeft1.trace";
file varLeft2trace : char_file open write_mode is "Top.MainvarLeft2.trace";
file varRighttrace : char_file open write_mode is "Top.MainvarRight.trace";
file varRight1trace : char_file open write_mode is "Top.MainvarRight1.trace";
file varRight2trace : char_file open write_mode is "Top.MainvarRight2.trace";
signal h0s_cond_synchscl000006d : std_logic_vector (0 downto 0);
signal h1s_cond_synchscl000006e : std_logic_vector (0 downto 0);
signal h1_cond1sT_synchscl000006f : std_logic_vector (0 downto 0);
signal h1_qssumsqssT_synchscl000006g :  std_logic_vector (48-1 downto 0);
signal h1_qssumssT_synchscl000006h :  std_logic_vector (48-1 downto 0);
signal h1_varLsT_synchscl000006i :  std_logic_vector (64-1 downto 0);
signal h1_condsT_synchscl000006j : std_logic_vector (0 downto 0);
signal h1sT_cond_synchscl000006k : std_logic_vector (0 downto 0);
signal h1sT_cond_sync1hscl000006l : std_logic_vector (0 downto 0);
signal h1sTE_cond_synchscl000006m : std_logic_vector (0 downto 0);
signal h1sTET_cond_synchscl000006n : std_logic_vector (0 downto 0);
signal h2s_cond_synchscl000006o : std_logic_vector (0 downto 0);
signal h2sE_cond_synchscl000006p : std_logic_vector (0 downto 0);
signal h3s_cond_synchscl000006q : std_logic_vector (0 downto 0);
signal h3sE_cond_synchscl000006r : std_logic_vector (0 downto 0);
signal h4s_cond_synchscl000006s : std_logic_vector (0 downto 0);
signal h5s_cond_synchscl000006t : std_logic_vector (0 downto 0);
signal h5sT_cond_synchscl000006u : std_logic_vector (0 downto 0);
signal h5sTT_cond_synchscl000006v : std_logic_vector (0 downto 0);
signal h5sTTT_cond_synchscl000006w : std_logic_vector (0 downto 0);
signal h5sTTT_cond_sync1hscl000006x : std_logic_vector (0 downto 0);
signal h5_condsTTE_synchscl000006y : std_logic_vector (0 downto 0);
signal h5sTTE_cond_synchscl000006z : std_logic_vector (0 downto 0);
signal h5sTTE_cond_sync1hscl0000070 : std_logic_vector (0 downto 0);
signal h5sTTEE_cond_synchscl0000071 : std_logic_vector (0 downto 0);
signal h6s_cond_synchscl0000072 : std_logic_vector (0 downto 0);
signal h7s_cond_synchscl0000073 : std_logic_vector (0 downto 0);
signal h7sT_cond_synchscl0000074 : std_logic_vector (0 downto 0);
signal h7_subsumsqssTT_synchscl0000075 :  std_logic_vector (48-1 downto 0);
signal h7_qssubsumssTT_synchscl0000076 :  std_logic_vector (48-1 downto 0);
signal h7_varRsTT_synchscl0000077 :  std_logic_vector (64-1 downto 0);
signal h7sTT_cond_synchscl0000078 : std_logic_vector (0 downto 0);
signal h7sT_cond_sync1hscl0000079 : std_logic_vector (0 downto 0);
signal h8_outpVars_rdys_synchscl000007a : std_logic_vector (0 downto 0);
signal h8_outp1_rdys_synchscl000007b : std_logic_vector (0 downto 0);
signal h8_outp_rdys_synchscl000007c : std_logic_vector (0 downto 0);
signal h8_h1s_finish4_rdys_synchscl000007d : std_logic_vector (0 downto 0);
signal h8_handlerForVarRCut_rdys_synchscl000007e : std_logic_vector (0 downto 0);
signal h8_h0_rdys_synchscl000007f : std_logic_vector (0 downto 0);
signal h8_h4_then_rdys_synchscl000007g : std_logic_vector (0 downto 0);
signal h8_h1sT_finish4_rdys_synchscl000007h : std_logic_vector (0 downto 0);
signal h8_h4_rdys_synchscl000007i : std_logic_vector (0 downto 0);
signal h8_h3_then_rdys_synchscl000007j : std_logic_vector (0 downto 0);
signal h8_h3_else_then_rdys_synchscl000007k : std_logic_vector (0 downto 0);
signal h8_h1sT_finish_rdys_synchscl000007l : std_logic_vector (0 downto 0);
signal h8_h3_else_rdys_synchscl000007m : std_logic_vector (0 downto 0);
signal h8_h1sTT_finish4_rdys_synchscl000007n : std_logic_vector (0 downto 0);
signal h8_h3_rdys_synchscl000007o : std_logic_vector (0 downto 0);
signal h8_h2_then_rdys_synchscl000007p : std_logic_vector (0 downto 0);
signal h8_h2_else_then_rdys_synchscl000007q : std_logic_vector (0 downto 0);
signal h8_h1sTTE_finish4_rdys_synchscl000007r : std_logic_vector (0 downto 0);
signal h8_h2_else_rdys_synchscl000007s : std_logic_vector (0 downto 0);
signal h8_h1sTT_finish_rdys_synchscl000007t : std_logic_vector (0 downto 0);
signal h8_h2_rdys_synchscl000007u : std_logic_vector (0 downto 0);
signal h8_h1_then_r_rdys_synchscl000007v : std_logic_vector (0 downto 0);
signal h8_h1_then_leftHappenings_synchscl000007w : std_logic_vector (0 downto 0);
signal h8_h1_then_enableRights_synchscl000007x : std_logic_vector (0 downto 0);
signal h8_h1_then_rdys_synchscl000007y : std_logic_vector (0 downto 0);
signal h8_h1sTTE_finish2_rdys_synchscl000007z : std_logic_vector (0 downto 0);
signal h8_h1_rdys_synchscl0000080 : std_logic_vector (0 downto 0);
signal h8_h5_then_then_then_r_rdys_synchscl0000081 : std_logic_vector (0 downto 0);
signal h8_h5_then_then_then_leftHappenings_synchscl0000082 : std_logic_vector (0 downto 0);
signal h8_h5_then_then_then_enableRights_synchscl0000083 : std_logic_vector (0 downto 0);
signal h8_h5_then_then_then_rdys_synchscl0000084 : std_logic_vector (0 downto 0);
signal h8_h5_then_then_else_r_rdys_synchscl0000085 : std_logic_vector (0 downto 0);
signal h8_h5_then_then_else_leftHappenings_synchscl0000086 : std_logic_vector (0 downto 0);
signal h8_h5_then_then_else_enableRights_synchscl0000087 : std_logic_vector (0 downto 0);
signal h8_h5_then_then_else_rdys_synchscl0000088 : std_logic_vector (0 downto 0);
signal h8_h5_then_then_rdys_synchscl0000089 : std_logic_vector (0 downto 0);
signal h8_h5_then_else_rdys_synchscl000008a : std_logic_vector (0 downto 0);
signal h8_h5_then_rdys_synchscl000008b : std_logic_vector (0 downto 0);
signal h8_inp_rdys_synchscl000008c : std_logic_vector (0 downto 0);
signal h8_h5_rdys_synchscl000008d : std_logic_vector (0 downto 0);
signal h8s_cond_synchscl000008e : std_logic_vector (0 downto 0);
signal h8s_cond_sync1hscl000008f : std_logic_vector (0 downto 0);
signal h8s_cond_sync2hscl000008g : std_logic_vector (0 downto 0);
signal h8s_cond_sync3hscl000008h : std_logic_vector (0 downto 0);
signal h8s_cond_sync4hscl000008i : std_logic_vector (0 downto 0);
signal h8s_cond_sync5hscl000008j : std_logic_vector (0 downto 0);
signal h8s_cond_sync6hscl000008k : std_logic_vector (0 downto 0);
signal h8s_cond_sync7hscl000008l : std_logic_vector (0 downto 0);
signal h8s_cond_sync8hscl000008m : std_logic_vector (0 downto 0);
signal h8s_cond_sync9hscl000008n : std_logic_vector (0 downto 0);
signal h8s_cond_sync10hscl000008o : std_logic_vector (0 downto 0);
signal h8s_cond_sync11hscl000008p : std_logic_vector (0 downto 0);

begin
i_TopMainhandlerForVar : entity work.proc_TopRdyCutStp0Isuint10 port map 
(rst => rst, clk => clk, reset_rdy_ena => reset_rdy_ena, outp_data => handlerForVarRCuthscl000001h_data, outp_ena => handlerForVarRCuthscl000001h_ena, inp_rdy_ena => handlerForVar_rdyhscl000001g_ena, reset_ena => reset_ena, inp_data => handlerForVarhscl000001f_data, inp_ena => handlerForVarhscl000001f_ena, outp_rdy_ena => handlerForVarRCut_rdyhscl000001e_ena)
;i_TopMainLInserter_h1sTTE1 : entity work.proc_TopLInserterStp0Isint16 port map 
 (rst => rst, clk => clk, outp_data => h1sTTE_finish4hscl000001d_data, outp_ena => h1sTTE_finish4hscl000001d_ena, inp_rdy_ena => h1sTTE_finish3_rdyhscl000001c_ena, reset_rdy_ena => reset_rdy_ena, reset_ena => reset_ena, inp_data => h1sTTE_finish3hscl000001b_data, inp_ena => h1sTTE_finish3hscl000001b_ena, outp_rdy_ena => h1sTTE_finish4_rdyhscl000001a_ena)
 ;i_TopMainPipe_h1sTTE0 : entity work.proc_TopPipeStp0Isint16 port map 
  (rst => rst, clk => clk, reset_rdy_ena => reset_rdy_ena, outp_data => h1sTTE_finish2hscl0000019_data, outp_ena => h1sTTE_finish2hscl0000019_ena, inp_rdy_ena => h1sTTE_finish1_rdyhscl0000012_ena, oBufFull_ena => Pipe_h1sTTE0BufFullhscl0000018_ena, reset_ena => reset_ena, inp_data => h1sTTE_finish1hscl0000015_data, inp_ena => h1sTTE_finish1hscl0000015_ena, outp_rdy_ena => h1sTTE_finish2_rdyhscl0000017_ena, oBufFull_rdy_ena => Pipe_h1sTTE0BufFull_rdyhscl0000016_ena)
  ;i_TopMainLInserter_h1sTTE0 : entity work.proc_TopLInserterStp0Isint16 port map 
   (rst => rst, clk => clk, outp_data => h1sTTE_finish1hscl0000015_data, outp_ena => h1sTTE_finish1hscl0000015_ena, inp_rdy_ena => h1sTTE_finish_rdyhscl0000014_ena, reset_rdy_ena => reset_rdy_ena, reset_ena => reset_ena, inp_data => h1sTTE_finishhscl0000013_data, inp_ena => h1sTTE_finishhscl0000013_ena, outp_rdy_ena => h1sTTE_finish1_rdyhscl0000012_ena)
   ;process (clk, rst) is
    variable defiPrintVar : std_logic_vector (0 downto 0) ;
    variable deficonflictCounter : integer ;
    variable endofoutpPrintVar : std_logic_vector (0 downto 0) ;
    variable endofoutpconflictCounter : integer ;
    variable endofoutp1PrintVar : std_logic_vector (0 downto 0) ;
    variable endofoutp1conflictCounter : integer ;
    variable h0_elseTransactionPrintVar : std_logic_vector (0 downto 0) ;
    variable h0_elseTransactionconflictCounter : integer ;
    variable h1_elseTransactionPrintVar : std_logic_vector (0 downto 0) ;
    variable h1_elseTransactionconflictCounter : integer ;
    variable h1_then_l_elseTransactionPrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h1_then_l_elseTransactionconflictCounter : integer ;
    variable h1_then_l_then_lastHappened0PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h1_then_l_then_lastHappened0conflictCounter : integer ;
    variable h1_then_l_then_lastHappened1PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h1_then_l_then_lastHappened1conflictCounter : integer ;
    variable h1_then_l_then_lastHappened2PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h1_then_l_then_lastHappened2conflictCounter : integer ;
    variable h1_then_l_then_p2_elseTransactionPrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h1_then_l_then_p2_elseTransactionconflictCounter : integer ;
    variable h1_then_leftHappenedPrintVar : std_logic_vector (0 downto 0) ;
    variable h1_then_leftHappenedconflictCounter : integer ;
    variable h2_elseTransactionPrintVar : std_logic_vector (0 downto 0) ;
    variable h2_elseTransactionconflictCounter : integer ;
    variable h2_else_elseTransactionPrintVar : std_logic_vector (0 downto 0) 
    ;
    variable h2_else_elseTransactionconflictCounter : integer ;
    variable h3_elseTransactionPrintVar : std_logic_vector (0 downto 0) ;
    variable h3_elseTransactionconflictCounter : integer ;
    variable h3_else_elseTransactionPrintVar : std_logic_vector (0 downto 0) 
    ;
    variable h3_else_elseTransactionconflictCounter : integer ;
    variable h4_elseTransactionPrintVar : std_logic_vector (0 downto 0) ;
    variable h4_elseTransactionconflictCounter : integer ;
    variable h5_elseTransactionPrintVar : std_logic_vector (0 downto 0) ;
    variable h5_elseTransactionconflictCounter : integer ;
    variable h5_then_elseTransactionPrintVar : std_logic_vector (0 downto 0) 
    ;
    variable h5_then_elseTransactionconflictCounter : integer ;
    variable h5_then_then_elseTransactionPrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h5_then_then_elseTransactionconflictCounter : integer ;
    variable h5_then_then_else_l_lastHappened0PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h5_then_then_else_l_lastHappened0conflictCounter : integer ;
    variable h5_then_then_else_l_lastHappened1PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h5_then_then_else_l_lastHappened1conflictCounter : integer ;
    variable h5_then_then_else_l_lastHappened2PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h5_then_then_else_l_lastHappened2conflictCounter : integer ;
    variable h5_then_then_else_l_p0_elseTransactionPrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h5_then_then_else_l_p0_elseTransactionconflictCounter : integer 
    ;
    variable h5_then_then_else_leftHappenedPrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h5_then_then_else_leftHappenedconflictCounter : integer ;
    variable h5_then_then_then_l_lastHappened0PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h5_then_then_then_l_lastHappened0conflictCounter : integer ;
    variable h5_then_then_then_l_lastHappened1PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h5_then_then_then_l_lastHappened1conflictCounter : integer ;
    variable h5_then_then_then_l_lastHappened2PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h5_then_then_then_l_lastHappened2conflictCounter : integer ;
    variable h5_then_then_then_leftHappenedPrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h5_then_then_then_leftHappenedconflictCounter : integer ;
    variable h6_elseTransactionPrintVar : std_logic_vector (0 downto 0) ;
    variable h6_elseTransactionconflictCounter : integer ;
    variable h7_elseTransactionPrintVar : std_logic_vector (0 downto 0) ;
    variable h7_elseTransactionconflictCounter : integer ;
    variable h7_then_lastHappened0PrintVar : std_logic_vector (0 downto 0) ;
    variable h7_then_lastHappened0conflictCounter : integer ;
    variable h7_then_lastHappened1PrintVar : std_logic_vector (0 downto 0) ;
    variable h7_then_lastHappened1conflictCounter : integer ;
    variable h7_then_p0_elseTransactionPrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p0_elseTransactionconflictCounter : integer ;
    variable h7_then_p0_then_lastHappened0PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p0_then_lastHappened0conflictCounter : integer ;
    variable h7_then_p0_then_lastHappened1PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p0_then_lastHappened1conflictCounter : integer ;
    variable h7_then_p0_then_lastHappened2PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p0_then_lastHappened2conflictCounter : integer ;
    variable h7_then_p0_then_p2_lastHappened0PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p0_then_p2_lastHappened0conflictCounter : integer ;
    variable h7_then_p0_then_p2_lastHappened1PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p0_then_p2_lastHappened1conflictCounter : integer ;
    variable h7_then_p0_then_p2_lastHappened2PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p0_then_p2_lastHappened2conflictCounter : integer ;
    variable h7_then_p0_then_p2_p2_elseTransactionPrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p0_then_p2_p2_elseTransactionconflictCounter : integer ;
    variable h7_then_p1_elseTransactionPrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_elseTransactionconflictCounter : integer ;
    variable h7_then_p1_then_lastHappened0PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened0conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened1PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened1conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened10PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened10conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened11PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened11conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened12PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened12conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened13PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened13conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened14PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened14conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened15PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened15conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened16PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened16conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened17PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened17conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened18PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened18conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened19PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened19conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened2PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened2conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened20PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened20conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened21PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened21conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened22PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened22conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened23PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened23conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened24PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened24conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened25PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened25conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened26PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened26conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened27PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened27conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened28PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened28conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened29PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened29conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened3PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened3conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened30PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened30conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened31PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened31conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened32PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened32conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened33PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened33conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened34PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened34conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened35PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened35conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened36PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened36conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened37PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened37conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened38PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened38conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened39PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened39conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened4PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened4conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened40PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened40conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened41PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened41conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened42PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened42conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened43PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened43conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened44PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened44conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened45PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened45conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened46PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened46conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened47PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened47conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened48PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened48conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened49PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened49conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened5PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened5conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened50PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened50conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened51PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened51conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened52PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened52conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened53PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened53conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened54PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened54conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened55PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened55conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened56PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened56conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened57PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened57conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened58PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened58conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened59PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened59conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened6PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened6conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened60PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened60conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened61PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened61conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened62PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened62conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened63PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened63conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened64PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened64conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened7PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened7conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened8PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened8conflictCounter : integer ;
    variable h7_then_p1_then_lastHappened9PrintVar : 
    std_logic_vector (0 downto 0) ;
    variable h7_then_p1_then_lastHappened9conflictCounter : integer ;
    variable iPrintVar :  std_logic_vector (10-1 downto 0) ;
    variable iconflictCounter : integer ;
    variable icoefmultPrintVar : arrticoefmult1(0 to 63) ;
    variable icoefmultconflictCounter : integer ;
    variable sumsPrintVar : arrtsums1(0 to 63) ;
    variable sumsconflictCounter : integer ;
    variable sumsqsPrintVar : arrtsumsqs1(0 to 63) ;
    variable sumsqsconflictCounter : integer ;
    variable varLeftPrintVar : arrtvarLeft1(0 to 63) ;
    variable varLeftconflictCounter : integer ;
    variable varLeft1PrintVar : arrtvarLeft11(0 to 63) ;
    variable varLeft1conflictCounter : integer ;
    variable varLeft2PrintVar : arrtvarLeft11(0 to 63) ;
    variable varLeft2conflictCounter : integer ;
    variable varRightPrintVar : arrtvarLeft1(0 to 63) ;
    variable varRightconflictCounter : integer ;
    variable varRight1PrintVar : arrtvarRight11(0 to 63) ;
    variable varRight1conflictCounter : integer ;
    variable varRight2PrintVar : arrtvarRight11(0 to 63) ;
    variable varRight2conflictCounter : integer ;
    variable rhs :  std_logic_vector (64-1 downto 0) ;
    variable rhs1 :  std_logic_vector (32-1 downto 0) ;
    variable rhs2 :  std_logic_vector (24-1 downto 0) ;
    variable tmp :  std_logic_vector (32-1 downto 0) ;
    variable rhs3 :  std_logic_vector (32-1 downto 0) ;
    variable tmp3 :  std_logic_vector (24-1 downto 0) ;
    variable rhs4 :  std_logic_vector (24-1 downto 0) ;
    variable rhs5 :  std_logic_vector (64-1 downto 0) ;
    variable rhs6 :  std_logic_vector (13-1 downto 0) ;
    variable rhs7 :  std_logic_vector (13-1 downto 0) ;
    variable rhs8 :  std_logic_vector (13-1 downto 0) ;
    variable rhs9 :  std_logic_vector (13-1 downto 0) ;
    variable rhs10 :  std_logic_vector (13-1 downto 0) ;
    variable rhs11 :  std_logic_vector (13-1 downto 0) ;
    variable rhs12 :  std_logic_vector (13-1 downto 0) ;
    variable rhs13 :  std_logic_vector (13-1 downto 0) ;
    variable rhs14 :  std_logic_vector (13-1 downto 0) ;
    variable rhs15 :  std_logic_vector (13-1 downto 0) ;
    variable rhs16 :  std_logic_vector (13-1 downto 0) ;
    variable rhs17 :  std_logic_vector (13-1 downto 0) ;
    variable rhs18 :  std_logic_vector (13-1 downto 0) ;
    variable rhs19 :  std_logic_vector (13-1 downto 0) ;
    variable rhs20 :  std_logic_vector (13-1 downto 0) ;
    variable rhs21 :  std_logic_vector (13-1 downto 0) ;
    variable rhs22 :  std_logic_vector (13-1 downto 0) ;
    variable rhs23 :  std_logic_vector (13-1 downto 0) ;
    variable rhs24 :  std_logic_vector (13-1 downto 0) ;
    variable rhs25 :  std_logic_vector (13-1 downto 0) ;
    variable rhs26 :  std_logic_vector (13-1 downto 0) ;
    variable rhs27 :  std_logic_vector (13-1 downto 0) ;
    variable rhs28 :  std_logic_vector (13-1 downto 0) ;
    variable rhs29 :  std_logic_vector (13-1 downto 0) ;
    variable rhs30 :  std_logic_vector (13-1 downto 0) ;
    variable rhs31 :  std_logic_vector (13-1 downto 0) ;
    variable rhs32 :  std_logic_vector (13-1 downto 0) ;
    variable rhs33 :  std_logic_vector (13-1 downto 0) ;
    variable rhs34 :  std_logic_vector (13-1 downto 0) ;
    variable rhs35 :  std_logic_vector (13-1 downto 0) ;
    variable rhs36 :  std_logic_vector (13-1 downto 0) ;
    variable rhs37 :  std_logic_vector (13-1 downto 0) ;
    variable rhs38 :  std_logic_vector (13-1 downto 0) ;
    variable rhs39 :  std_logic_vector (13-1 downto 0) ;
    variable rhs40 :  std_logic_vector (13-1 downto 0) ;
    variable rhs41 :  std_logic_vector (13-1 downto 0) ;
    variable rhs42 :  std_logic_vector (13-1 downto 0) ;
    variable rhs43 :  std_logic_vector (13-1 downto 0) ;
    variable rhs44 :  std_logic_vector (13-1 downto 0) ;
    variable rhs45 :  std_logic_vector (13-1 downto 0) ;
    variable rhs46 :  std_logic_vector (13-1 downto 0) ;
    variable rhs47 :  std_logic_vector (13-1 downto 0) ;
    variable rhs48 :  std_logic_vector (13-1 downto 0) ;
    variable rhs49 :  std_logic_vector (13-1 downto 0) ;
    variable rhs50 :  std_logic_vector (13-1 downto 0) ;
    variable rhs51 :  std_logic_vector (13-1 downto 0) ;
    variable rhs52 :  std_logic_vector (13-1 downto 0) ;
    variable rhs53 :  std_logic_vector (13-1 downto 0) ;
    variable rhs54 :  std_logic_vector (13-1 downto 0) ;
    variable rhs55 :  std_logic_vector (13-1 downto 0) ;
    variable rhs56 :  std_logic_vector (13-1 downto 0) ;
    variable rhs57 :  std_logic_vector (13-1 downto 0) ;
    variable rhs58 :  std_logic_vector (13-1 downto 0) ;
    variable rhs59 :  std_logic_vector (13-1 downto 0) ;
    variable rhs60 :  std_logic_vector (13-1 downto 0) ;
    variable rhs61 :  std_logic_vector (13-1 downto 0) ;
    variable rhs62 :  std_logic_vector (13-1 downto 0) ;
    variable rhs63 :  std_logic_vector (13-1 downto 0) ;
    variable rhs64 :  std_logic_vector (13-1 downto 0) ;
    variable rhs65 :  std_logic_vector (13-1 downto 0) ;
    variable rhs66 :  std_logic_vector (13-1 downto 0) ;
    variable rhs67 :  std_logic_vector (13-1 downto 0) ;
    variable rhs68 :  std_logic_vector (13-1 downto 0) ;
    variable rhs69 :  std_logic_vector (13-1 downto 0) ;
    variable tmp69 : std_logic_vector (0 downto 0) ;
    variable tmp70 : std_logic_vector (0 downto 0) ;
    variable tmp71 : std_logic_vector (0 downto 0) ;
    variable tmp72 : std_logic_vector (0 downto 0) ;
    variable tmp73 : std_logic_vector (0 downto 0) ;
    variable tmp74 : std_logic_vector (0 downto 0) ;
    variable tmp75 : std_logic_vector (0 downto 0) ;
    variable tmp76 : std_logic_vector (0 downto 0) ;
    variable tmp77 : std_logic_vector (0 downto 0) ;
    variable tmp78 : std_logic_vector (0 downto 0) ;
    variable tmp79 : std_logic_vector (0 downto 0) ;
    variable tmp80 : std_logic_vector (0 downto 0) ;
    begin
      if clk'event and clk = '1' then
        deficonflictCounter := 0 ;
        endofoutpconflictCounter := 0 ;
        endofoutp1conflictCounter := 0 ;
        h0_elseTransactionconflictCounter := 0 ;
        h1_elseTransactionconflictCounter := 0 ;
        h1_then_l_elseTransactionconflictCounter := 0 ;
        h1_then_l_then_lastHappened0conflictCounter := 0 ;
        h1_then_l_then_lastHappened1conflictCounter := 0 ;
        h1_then_l_then_lastHappened2conflictCounter := 0 ;
        h1_then_l_then_p2_elseTransactionconflictCounter := 0 ;
        h1_then_leftHappenedconflictCounter := 0 ;
        h2_elseTransactionconflictCounter := 0 ;
        h2_else_elseTransactionconflictCounter := 0 ;
        h3_elseTransactionconflictCounter := 0 ;
        h3_else_elseTransactionconflictCounter := 0 ;
        h4_elseTransactionconflictCounter := 0 ;
        h5_elseTransactionconflictCounter := 0 ;
        h5_then_elseTransactionconflictCounter := 0 ;
        h5_then_then_elseTransactionconflictCounter := 0 ;
        h5_then_then_else_l_lastHappened0conflictCounter := 0 ;
        h5_then_then_else_l_lastHappened1conflictCounter := 0 ;
        h5_then_then_else_l_lastHappened2conflictCounter := 0 ;
        h5_then_then_else_l_p0_elseTransactionconflictCounter := 0 ;
        h5_then_then_else_leftHappenedconflictCounter := 0 ;
        h5_then_then_then_l_lastHappened0conflictCounter := 0 ;
        h5_then_then_then_l_lastHappened1conflictCounter := 0 ;
        h5_then_then_then_l_lastHappened2conflictCounter := 0 ;
        h5_then_then_then_leftHappenedconflictCounter := 0 ;
        h6_elseTransactionconflictCounter := 0 ;
        h7_elseTransactionconflictCounter := 0 ;
        h7_then_lastHappened0conflictCounter := 0 ;
        h7_then_lastHappened1conflictCounter := 0 ;
        h7_then_p0_elseTransactionconflictCounter := 0 ;
        h7_then_p0_then_lastHappened0conflictCounter := 0 ;
        h7_then_p0_then_lastHappened1conflictCounter := 0 ;
        h7_then_p0_then_lastHappened2conflictCounter := 0 ;
        h7_then_p0_then_p2_lastHappened0conflictCounter := 0 ;
        h7_then_p0_then_p2_lastHappened1conflictCounter := 0 ;
        h7_then_p0_then_p2_lastHappened2conflictCounter := 0 ;
        h7_then_p0_then_p2_p2_elseTransactionconflictCounter := 0 ;
        h7_then_p1_elseTransactionconflictCounter := 0 ;
        h7_then_p1_then_lastHappened0conflictCounter := 0 ;
        h7_then_p1_then_lastHappened1conflictCounter := 0 ;
        h7_then_p1_then_lastHappened10conflictCounter := 0 ;
        h7_then_p1_then_lastHappened11conflictCounter := 0 ;
        h7_then_p1_then_lastHappened12conflictCounter := 0 ;
        h7_then_p1_then_lastHappened13conflictCounter := 0 ;
        h7_then_p1_then_lastHappened14conflictCounter := 0 ;
        h7_then_p1_then_lastHappened15conflictCounter := 0 ;
        h7_then_p1_then_lastHappened16conflictCounter := 0 ;
        h7_then_p1_then_lastHappened17conflictCounter := 0 ;
        h7_then_p1_then_lastHappened18conflictCounter := 0 ;
        h7_then_p1_then_lastHappened19conflictCounter := 0 ;
        h7_then_p1_then_lastHappened2conflictCounter := 0 ;
        h7_then_p1_then_lastHappened20conflictCounter := 0 ;
        h7_then_p1_then_lastHappened21conflictCounter := 0 ;
        h7_then_p1_then_lastHappened22conflictCounter := 0 ;
        h7_then_p1_then_lastHappened23conflictCounter := 0 ;
        h7_then_p1_then_lastHappened24conflictCounter := 0 ;
        h7_then_p1_then_lastHappened25conflictCounter := 0 ;
        h7_then_p1_then_lastHappened26conflictCounter := 0 ;
        h7_then_p1_then_lastHappened27conflictCounter := 0 ;
        h7_then_p1_then_lastHappened28conflictCounter := 0 ;
        h7_then_p1_then_lastHappened29conflictCounter := 0 ;
        h7_then_p1_then_lastHappened3conflictCounter := 0 ;
        h7_then_p1_then_lastHappened30conflictCounter := 0 ;
        h7_then_p1_then_lastHappened31conflictCounter := 0 ;
        h7_then_p1_then_lastHappened32conflictCounter := 0 ;
        h7_then_p1_then_lastHappened33conflictCounter := 0 ;
        h7_then_p1_then_lastHappened34conflictCounter := 0 ;
        h7_then_p1_then_lastHappened35conflictCounter := 0 ;
        h7_then_p1_then_lastHappened36conflictCounter := 0 ;
        h7_then_p1_then_lastHappened37conflictCounter := 0 ;
        h7_then_p1_then_lastHappened38conflictCounter := 0 ;
        h7_then_p1_then_lastHappened39conflictCounter := 0 ;
        h7_then_p1_then_lastHappened4conflictCounter := 0 ;
        h7_then_p1_then_lastHappened40conflictCounter := 0 ;
        h7_then_p1_then_lastHappened41conflictCounter := 0 ;
        h7_then_p1_then_lastHappened42conflictCounter := 0 ;
        h7_then_p1_then_lastHappened43conflictCounter := 0 ;
        h7_then_p1_then_lastHappened44conflictCounter := 0 ;
        h7_then_p1_then_lastHappened45conflictCounter := 0 ;
        h7_then_p1_then_lastHappened46conflictCounter := 0 ;
        h7_then_p1_then_lastHappened47conflictCounter := 0 ;
        h7_then_p1_then_lastHappened48conflictCounter := 0 ;
        h7_then_p1_then_lastHappened49conflictCounter := 0 ;
        h7_then_p1_then_lastHappened5conflictCounter := 0 ;
        h7_then_p1_then_lastHappened50conflictCounter := 0 ;
        h7_then_p1_then_lastHappened51conflictCounter := 0 ;
        h7_then_p1_then_lastHappened52conflictCounter := 0 ;
        h7_then_p1_then_lastHappened53conflictCounter := 0 ;
        h7_then_p1_then_lastHappened54conflictCounter := 0 ;
        h7_then_p1_then_lastHappened55conflictCounter := 0 ;
        h7_then_p1_then_lastHappened56conflictCounter := 0 ;
        h7_then_p1_then_lastHappened57conflictCounter := 0 ;
        h7_then_p1_then_lastHappened58conflictCounter := 0 ;
        h7_then_p1_then_lastHappened59conflictCounter := 0 ;
        h7_then_p1_then_lastHappened6conflictCounter := 0 ;
        h7_then_p1_then_lastHappened60conflictCounter := 0 ;
        h7_then_p1_then_lastHappened61conflictCounter := 0 ;
        h7_then_p1_then_lastHappened62conflictCounter := 0 ;
        h7_then_p1_then_lastHappened63conflictCounter := 0 ;
        h7_then_p1_then_lastHappened64conflictCounter := 0 ;
        h7_then_p1_then_lastHappened7conflictCounter := 0 ;
        h7_then_p1_then_lastHappened8conflictCounter := 0 ;
        h7_then_p1_then_lastHappened9conflictCounter := 0 ;
        iconflictCounter := 0 ;
        icoefmultconflictCounter := 0 ;
        sumsconflictCounter := 0 ;
        sumsqsconflictCounter := 0 ;
        varLeftconflictCounter := 0 ;
        varLeft1conflictCounter := 0 ;
        varLeft2conflictCounter := 0 ;
        varRightconflictCounter := 0 ;
        varRight1conflictCounter := 0 ;
        varRight2conflictCounter := 0 ;
        rhs := h1_varLsT_synchscl000006i ;
        if h1s_cond_synchscl000006e(0)='1' then
          if h1sT_cond_sync1hscl000006l(0)='1' then
            null;
          else
            if h1sTE_cond_synchscl000006m(0)='1' then
              if h1sTET_cond_synchscl000006n(0)='1' then
                endofoutpPrintVar := endofoutphscl0000036 ;
                fprint_stringPtr(endofoutptrace,   toStringUnsigned(endofoutpPrintVar));
                fprint_string(endofoutptrace,  newline);
                endofoutpconflictCounter := endofoutpconflictCounter + 1;
                assert endofoutpconflictCounter <= 1 report "conflict when writing endofoutp" severity failure ; 
                endofoutphscl0000036 <= 
                 conv_std_logic_vector(std_logic_vector'(B"1")) ;
              else
                null;
              end if;
              varLefthscl0000067(notCheck(0 +  conv_integer_bound_unsigned
                                              (conv_std_logic_vector(conv_std_logic_vector
                                                                    (bc_unsigned_sub
                                                                    (ihscl0000063,   conv_std_logic_vector
                                                                    (1,  10)))),  0),  0,  63)) <= rhs;
            else
              null;
            end if;
          end if;
        else
          null;
        end if;
        rhs1 := 
        conv_std_logic_vector(conv_std_logic_vector(bc_signed_emul(inp_data.p0,  inp_data.p0))) 
        ;
        rhs2 := bc_signed_c_sxt(inp_data.p0,  24) ;
        tmp := 
        arrayTrim(sumsqshscl0000066,  conv_std_logic_vector(conv_std_logic_vector
                                                            (bc_unsigned_sub
                                                             (ihscl0000063,   conv_std_logic_vector
                                                                    (1,  10))))) 
        ;
        rhs3 := 
        bc_unsigned_add(tmp,  conv_std_logic_vector(conv_std_logic_vector
                                                    (bc_signed_emul(inp_data.p0,  inp_data.p0)))) 
        ;
        tmp3 := 
        arrayTrim(sumshscl0000065,  conv_std_logic_vector(conv_std_logic_vector
                                                          (bc_unsigned_sub
                                                           (ihscl0000063,   conv_std_logic_vector
                                                                    (1,  10))))) 
        ;
        rhs4 := bc_signed_add(tmp3,  bc_signed_c_sxt(inp_data.p0,  24)) ;
        if h5s_cond_synchscl000006t(0)='1' then
          if h5sT_cond_synchscl000006u(0)='1' then
            if h5sTT_cond_synchscl000006v(0)='1' then
              if h5sTTT_cond_sync1hscl000006x(0)='1' then
                null;
              else
                sumshscl0000065(notCheck(0 +  conv_integer_bound_unsigned
                                             (ihscl0000063,  0),  0,  63)) <= rhs2;
                sumsqshscl0000066(notCheck(0 +  conv_integer_bound_unsigned
                                               (ihscl0000063,  0),  0,  63)) <= rhs1;
                iPrintVar := ihscl0000063 ;
                fprint_stringPtr(itrace,   toStringUnsigned(iPrintVar));
                fprint_string(itrace,  newline);
                iconflictCounter := iconflictCounter + 1;
                assert iconflictCounter <= 1 report "conflict when writing i" severity failure ; 
                ihscl0000063 <= 
                bc_unsigned_add(ihscl0000063,   conv_std_logic_vector(1,  10)) 
                ;
              end if;
            else
              if h5sTTE_cond_sync1hscl0000070(0)='1' then
                null;
              else
                sumshscl0000065(notCheck(0 +  conv_integer_bound_unsigned
                                             (ihscl0000063,  0),  0,  63)) <= rhs4;
                sumsqshscl0000066(notCheck(0 +  conv_integer_bound_unsigned
                                               (ihscl0000063,  0),  0,  63)) <= rhs3;
                if h5sTTEE_cond_synchscl0000071(0)='1' then
                  iPrintVar := ihscl0000063 ;
                  fprint_stringPtr(itrace,   toStringUnsigned(iPrintVar));
                  fprint_string(itrace,  newline);
                  iconflictCounter := iconflictCounter + 1;
                  assert iconflictCounter <= 1 report "conflict when writing i" severity failure ; 
                  ihscl0000063 <= 
                  bc_unsigned_add(ihscl0000063,   conv_std_logic_vector
                                                 (2,  10)) ;
                else
                  iPrintVar := ihscl0000063 ;
                  fprint_stringPtr(itrace,   toStringUnsigned(iPrintVar));
                  fprint_string(itrace,  newline);
                  iconflictCounter := iconflictCounter + 1;
                  assert iconflictCounter <= 1 report "conflict when writing i" severity failure ; 
                  ihscl0000063 <= 
                  bc_unsigned_add(ihscl0000063,   conv_std_logic_vector
                                                 (1,  10)) ;
                end if;
              end if;
            end if;
          else
            null;
          end if;
        else
          null;
        end if;
        rhs5 := h7_varRsTT_synchscl0000077 ;
        rhs6 :=  conv_std_logic_vector(65,  13) ;
        rhs7 :=  conv_std_logic_vector(66,  13) ;
        rhs8 :=  conv_std_logic_vector(67,  13) ;
        rhs9 :=  conv_std_logic_vector(68,  13) ;
        rhs10 :=  conv_std_logic_vector(69,  13) ;
        rhs11 :=  conv_std_logic_vector(70,  13) ;
        rhs12 :=  conv_std_logic_vector(71,  13) ;
        rhs13 :=  conv_std_logic_vector(73,  13) ;
        rhs14 :=  conv_std_logic_vector(74,  13) ;
        rhs15 :=  conv_std_logic_vector(75,  13) ;
        rhs16 :=  conv_std_logic_vector(77,  13) ;
        rhs17 :=  conv_std_logic_vector(78,  13) ;
        rhs18 :=  conv_std_logic_vector(80,  13) ;
        rhs19 :=  conv_std_logic_vector(81,  13) ;
        rhs20 :=  conv_std_logic_vector(83,  13) ;
        rhs21 :=  conv_std_logic_vector(85,  13) ;
        rhs22 :=  conv_std_logic_vector(87,  13) ;
        rhs23 :=  conv_std_logic_vector(89,  13) ;
        rhs24 :=  conv_std_logic_vector(91,  13) ;
        rhs25 :=  conv_std_logic_vector(93,  13) ;
        rhs26 :=  conv_std_logic_vector(95,  13) ;
        rhs27 :=  conv_std_logic_vector(97,  13) ;
        rhs28 :=  conv_std_logic_vector(99,  13) ;
        rhs29 :=  conv_std_logic_vector(102,  13) ;
        rhs30 :=  conv_std_logic_vector(105,  13) ;
        rhs31 :=  conv_std_logic_vector(107,  13) ;
        rhs32 :=  conv_std_logic_vector(110,  13) ;
        rhs33 :=  conv_std_logic_vector(113,  13) ;
        rhs34 :=  conv_std_logic_vector(117,  13) ;
        rhs35 :=  conv_std_logic_vector(120,  13) ;
        rhs36 :=  conv_std_logic_vector(124,  13) ;
        rhs37 :=  conv_std_logic_vector(128,  13) ;
        rhs38 :=  conv_std_logic_vector(132,  13) ;
        rhs39 :=  conv_std_logic_vector(136,  13) ;
        rhs40 :=  conv_std_logic_vector(141,  13) ;
        rhs41 :=  conv_std_logic_vector(146,  13) ;
        rhs42 :=  conv_std_logic_vector(151,  13) ;
        rhs43 :=  conv_std_logic_vector(157,  13) ;
        rhs44 :=  conv_std_logic_vector(163,  13) ;
        rhs45 :=  conv_std_logic_vector(170,  13) ;
        rhs46 :=  conv_std_logic_vector(178,  13) ;
        rhs47 :=  conv_std_logic_vector(186,  13) ;
        rhs48 :=  conv_std_logic_vector(195,  13) ;
        rhs49 :=  conv_std_logic_vector(204,  13) ;
        rhs50 :=  conv_std_logic_vector(215,  13) ;
        rhs51 :=  conv_std_logic_vector(227,  13) ;
        rhs52 :=  conv_std_logic_vector(240,  13) ;
        rhs53 :=  conv_std_logic_vector(256,  13) ;
        rhs54 :=  conv_std_logic_vector(273,  13) ;
        rhs55 :=  conv_std_logic_vector(292,  13) ;
        rhs56 :=  conv_std_logic_vector(315,  13) ;
        rhs57 :=  conv_std_logic_vector(341,  13) ;
        rhs58 :=  conv_std_logic_vector(372,  13) ;
        rhs59 :=  conv_std_logic_vector(409,  13) ;
        rhs60 :=  conv_std_logic_vector(455,  13) ;
        rhs61 :=  conv_std_logic_vector(512,  13) ;
        rhs62 :=  conv_std_logic_vector(585,  13) ;
        rhs63 :=  conv_std_logic_vector(682,  13) ;
        rhs64 :=  conv_std_logic_vector(819,  13) ;
        rhs65 :=  conv_std_logic_vector(1024,  13) ;
        rhs66 :=  conv_std_logic_vector(1365,  13) ;
        rhs67 :=  conv_std_logic_vector(2048,  13) ;
        rhs68 :=  conv_std_logic_vector(4096,  13) ;
        rhs69 :=  conv_std_logic_vector(0,  13) ;
        if h7s_cond_synchscl0000073(0)='1' then
          if h7sT_cond_sync1hscl0000079(0)='1' then
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector(0,  10),  0),  0,  63)) <= rhs69;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector(1,  10),  0),  0,  63)) <= rhs68;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector(2,  10),  0),  0,  63)) <= rhs67;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector(3,  10),  0),  0,  63)) <= rhs66;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector(4,  10),  0),  0,  63)) <= rhs65;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector(5,  10),  0),  0,  63)) <= rhs64;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector(6,  10),  0),  0,  63)) <= rhs63;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector(7,  10),  0),  0,  63)) <= rhs62;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector(8,  10),  0),  0,  63)) <= rhs61;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector(9,  10),  0),  0,  63)) <= rhs60;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (10,  10),  0),  0,  63)) <= rhs59;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (11,  10),  0),  0,  63)) <= rhs58;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (12,  10),  0),  0,  63)) <= rhs57;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (13,  10),  0),  0,  63)) <= rhs56;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (14,  10),  0),  0,  63)) <= rhs55;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (15,  10),  0),  0,  63)) <= rhs54;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (16,  10),  0),  0,  63)) <= rhs53;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (17,  10),  0),  0,  63)) <= rhs52;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (18,  10),  0),  0,  63)) <= rhs51;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (19,  10),  0),  0,  63)) <= rhs50;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (20,  10),  0),  0,  63)) <= rhs49;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (21,  10),  0),  0,  63)) <= rhs48;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (22,  10),  0),  0,  63)) <= rhs47;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (23,  10),  0),  0,  63)) <= rhs46;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (24,  10),  0),  0,  63)) <= rhs45;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (25,  10),  0),  0,  63)) <= rhs44;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (26,  10),  0),  0,  63)) <= rhs43;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (27,  10),  0),  0,  63)) <= rhs42;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (28,  10),  0),  0,  63)) <= rhs41;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (29,  10),  0),  0,  63)) <= rhs40;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (30,  10),  0),  0,  63)) <= rhs39;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (31,  10),  0),  0,  63)) <= rhs38;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (32,  10),  0),  0,  63)) <= rhs37;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (33,  10),  0),  0,  63)) <= rhs36;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (34,  10),  0),  0,  63)) <= rhs35;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (35,  10),  0),  0,  63)) <= rhs34;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (36,  10),  0),  0,  63)) <= rhs33;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (37,  10),  0),  0,  63)) <= rhs32;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (38,  10),  0),  0,  63)) <= rhs31;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (39,  10),  0),  0,  63)) <= rhs30;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (40,  10),  0),  0,  63)) <= rhs29;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (41,  10),  0),  0,  63)) <= rhs28;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (42,  10),  0),  0,  63)) <= rhs27;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (43,  10),  0),  0,  63)) <= rhs26;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (44,  10),  0),  0,  63)) <= rhs25;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (45,  10),  0),  0,  63)) <= rhs24;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (46,  10),  0),  0,  63)) <= rhs23;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (47,  10),  0),  0,  63)) <= rhs22;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (48,  10),  0),  0,  63)) <= rhs21;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (49,  10),  0),  0,  63)) <= rhs20;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (50,  10),  0),  0,  63)) <= rhs19;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (51,  10),  0),  0,  63)) <= rhs18;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (52,  10),  0),  0,  63)) <= rhs17;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (53,  10),  0),  0,  63)) <= rhs16;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (54,  10),  0),  0,  63)) <= rhs15;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (55,  10),  0),  0,  63)) <= rhs14;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (56,  10),  0),  0,  63)) <= rhs13;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (57,  10),  0),  0,  63)) <= rhs12;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (58,  10),  0),  0,  63)) <= rhs11;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (59,  10),  0),  0,  63)) <= rhs10;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (60,  10),  0),  0,  63)) <= rhs9;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (61,  10),  0),  0,  63)) <= rhs8;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (62,  10),  0),  0,  63)) <= rhs7;
            icoefmulthscl0000064(notCheck(0 +  conv_integer_bound_unsigned
                                              ( conv_std_logic_vector
                                               (63,  10),  0),  0,  63)) <= rhs6;
            defiPrintVar := defihscl0000035 ;
            fprint_stringPtr(defitrace,  toString(defiPrintVar));
            fprint_string(defitrace,  newline);
            deficonflictCounter := deficonflictCounter + 1;
            assert deficonflictCounter <= 1 report "conflict when writing defi" severity failure ; 
            defihscl0000035 <= std_logic_vector'(B"0") ;
          else
            null;
          end if;
          if h7sT_cond_synchscl0000074(0)='1' then
            if h7sTT_cond_synchscl0000078(0)='1' then
              endofoutp1PrintVar := endofoutp1hscl0000037 ;
              fprint_stringPtr(endofoutp1trace,   toStringUnsigned(endofoutp1PrintVar));
              fprint_string(endofoutp1trace,  newline);
              endofoutp1conflictCounter := endofoutp1conflictCounter + 1;
              assert endofoutp1conflictCounter <= 1 report "conflict when writing endofoutp1" severity failure ; 
              endofoutp1hscl0000037 <= 
               conv_std_logic_vector(std_logic_vector'(B"1")) ;
            else
              null;
            end if;
            varRighthscl000006a(notCheck(0 +  conv_integer_bound_unsigned
                                             (conv_std_logic_vector(conv_std_logic_vector
                                                                    (bc_unsigned_sub
                                                                    (ihscl0000063,   conv_std_logic_vector
                                                                    (64,  10)))),  0),  0,  63)) <= rhs5;
            iPrintVar := ihscl0000063 ;
            fprint_stringPtr(itrace,   toStringUnsigned(iPrintVar));
            fprint_string(itrace,  newline);
            iconflictCounter := iconflictCounter + 1;
            assert iconflictCounter <= 1 report "conflict when writing i" severity failure ; 
            ihscl0000063 <= 
            bc_unsigned_add(ihscl0000063,   conv_std_logic_vector(1,  10)) ;
          else
            null;
          end if;
        else
          null;
        end if;
        if conv_boolean(h8_h5_then_then_else_rdys_synchscl0000088) then
          tmp69 := (0 => '0') ;
        else
          tmp69 := (0 => '1') ;
        end if;
        if conv_boolean((0 => h5_then_then_elseEnablehscl000002h_ena)) then
          tmp70 := tmp69 ;
        else
          tmp70 := h5_then_then_elseTransactionhscl000003n ;
        end if;
        if conv_boolean((0 => reset_ena)) then
          tmp71 := (0 => '0') ;
        else
          tmp71 := tmp70 ;
        end if;
        if conv_boolean(h8_h5_then_then_else_leftHappenings_synchscl0000086) then
          tmp72 := (0 => '1') ;
        else
          tmp72 := h5_then_then_else_leftHappenedhscl000003s ;
        end if;
        if conv_boolean(h8_h5_then_then_else_r_rdys_synchscl0000085) then
          tmp73 := (0 => '0') ;
        else
          tmp73 := tmp72 ;
        end if;
        if conv_boolean((0 => reset_ena)) then
          tmp74 := (0 => '0') ;
        else
          tmp74 := tmp73 ;
        end if;
        if conv_boolean(h8_h5_then_then_then_leftHappenings_synchscl0000082) then
          tmp75 := (0 => '1') ;
        else
          tmp75 := h5_then_then_then_leftHappenedhscl000003w ;
        end if;
        if conv_boolean(h8_h5_then_then_then_r_rdys_synchscl0000081) then
          tmp76 := (0 => '0') ;
        else
          tmp76 := tmp75 ;
        end if;
        if conv_boolean((0 => reset_ena)) then
          tmp77 := (0 => '0') ;
        else
          tmp77 := tmp76 ;
        end if;
        if conv_boolean(h8_h1_then_leftHappenings_synchscl000007w) then
          tmp78 := (0 => '1') ;
        else
          tmp78 := h1_then_leftHappenedhscl000003f ;
        end if;
        if conv_boolean(h8_h1_then_r_rdys_synchscl000007v) then
          tmp79 := (0 => '0') ;
        else
          tmp79 := tmp78 ;
        end if;
        if conv_boolean((0 => reset_ena)) then
          tmp80 := (0 => '0') ;
        else
          tmp80 := tmp79 ;
        end if;
        h1_then_leftHappenedPrintVar := h1_then_leftHappenedhscl000003f ;
        fprint_stringPtr(h1_then_leftHappenedtrace,  toString(h1_then_leftHappenedPrintVar));
        fprint_string(h1_then_leftHappenedtrace,  newline);
        h1_then_leftHappenedconflictCounter := h1_then_leftHappenedconflictCounter + 1;
        assert h1_then_leftHappenedconflictCounter <= 1 report "conflict when writing h1_then_leftHappened" severity failure ; 
        h1_then_leftHappenedhscl000003f <= tmp80 ;
        h5_then_then_then_leftHappenedPrintVar := 
        h5_then_then_then_leftHappenedhscl000003w ;
        fprint_stringPtr(h5_then_then_then_leftHappenedtrace,  toString
                                                               (h5_then_then_then_leftHappenedPrintVar));
        fprint_string(h5_then_then_then_leftHappenedtrace,  newline);
        h5_then_then_then_leftHappenedconflictCounter := h5_then_then_then_leftHappenedconflictCounter + 1;
        assert h5_then_then_then_leftHappenedconflictCounter <= 1 report "conflict when writing h5_then_then_then_leftHappened" severity failure ; 
        h5_then_then_then_leftHappenedhscl000003w <= tmp77 ;
        h5_then_then_else_leftHappenedPrintVar := 
        h5_then_then_else_leftHappenedhscl000003s ;
        fprint_stringPtr(h5_then_then_else_leftHappenedtrace,  toString
                                                               (h5_then_then_else_leftHappenedPrintVar));
        fprint_string(h5_then_then_else_leftHappenedtrace,  newline);
        h5_then_then_else_leftHappenedconflictCounter := h5_then_then_else_leftHappenedconflictCounter + 1;
        assert h5_then_then_else_leftHappenedconflictCounter <= 1 report "conflict when writing h5_then_then_else_leftHappened" severity failure ; 
        h5_then_then_else_leftHappenedhscl000003s <= tmp74 ;
        h5_then_then_elseTransactionPrintVar := 
        h5_then_then_elseTransactionhscl000003n ;
        fprint_stringPtr(h5_then_then_elseTransactiontrace,  toString
                                                             (h5_then_then_elseTransactionPrintVar));
        fprint_string(h5_then_then_elseTransactiontrace,  newline);
        h5_then_then_elseTransactionconflictCounter := h5_then_then_elseTransactionconflictCounter + 1;
        assert h5_then_then_elseTransactionconflictCounter <= 1 report "conflict when writing h5_then_then_elseTransaction" severity failure ; 
        h5_then_then_elseTransactionhscl000003n <= tmp71 ;
      end if;
    end process;
    process (reset_ena, handlerForVarRCuthscl000001h_data, handlerForVarRCuthscl000001h_ena) 
    is
    variable s_condExpr : std_logic_vector (0 downto 0) ;
    variable s_cond : std_logic ;
    variable h0s_cond_synchscl000006d_data_dummy : 
    std_logic_vector (0 downto 0) ;
    begin
      h0_thenEnablehscl000001j_ena <= '0' ;
      
      
      null;
      h0s_cond_synchscl000006d_data_dummy := 
      zero(h0s_cond_synchscl000006d_data_dummy) ;
      h0s_cond_synchscl000006d <= h0s_cond_synchscl000006d_data_dummy ;
      
      s_condExpr := 
      and2(not2((0 => '0')),  and2(not2((0 => reset_ena)),  (0 => '1'))) ;
      s_cond := (s_condExpr(0)) and handlerForVarRCuthscl000001h_ena ;
      h0s_cond_synchscl000006d <= (0 => s_cond) ;
      if (s_cond='1') then
        h0_thenEnablehscl000001j_ena <= '1' ;
        null;
      else
        null;
      end if;
      null;
    end process;
    process (sumshscl0000065, sumsqshscl0000066, icoefmulthscl0000064, h1sTTE_finish2hscl0000019_ena, h1_then_rightEnablehscl000001s_ena, endofoutphscl0000036, h1sTTE_finish2hscl0000019_data, ihscl0000063, h1_then_leftHappenedhscl000003f) 
    is
    variable s_condExpr : std_logic_vector (0 downto 0) ;
    variable s_cond : std_logic ;
    variable cond1_sT : std_logic_vector (0 downto 0) ;
    variable qssumsqs_sT :  std_logic_vector (48-1 downto 0) ;
    variable tmp :  std_logic_vector (32-1 downto 0) ;
    variable qssums_sT :  std_logic_vector (48-1 downto 0) ;
    variable tmp1 :  std_logic_vector (24-1 downto 0) ;
    variable tmp2 :  std_logic_vector (24-1 downto 0) ;
    variable varL_sT :  std_logic_vector (64-1 downto 0) ;
    variable tmp3 :  std_logic_vector (64-1 downto 0) ;
    variable tmp4 :  std_logic_vector (48-1 downto 0) ;
    variable tmp5 :  std_logic_vector (64-1 downto 0) ;
    variable cond_sT : std_logic_vector (0 downto 0) ;
    variable sT_condExpr : std_logic_vector (0 downto 0) ;
    variable sT_cond : std_logic ;
    variable sT_condExpr5 : std_logic_vector (0 downto 0) ;
    variable sT_cond5 : std_logic ;
    variable sTE_condExpr : std_logic_vector (0 downto 0) ;
    variable sTE_cond : std_logic ;
    variable sTET_condExpr : std_logic_vector (0 downto 0) ;
    variable sTET_cond : std_logic ;
    variable h1sT_cond_sync1hscl000006l_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h1s_cond_synchscl000006e_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h1sT_cond_synchscl000006k_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h1sTE_cond_synchscl000006m_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h1sTET_cond_synchscl000006n_data_dummy : 
    std_logic_vector (0 downto 0) ;
    begin
      h1_then_l_thenEnablehscl000001o_ena <= '0' ;
      h1_then_enablehscl000001m_ena <= '0' ;
      h1_thenEnablehscl000001l_ena <= '0' ;
      h1sTTE_finish3hscl000001b_ena <= '0' ;
      h1_then_l_then_p2_thenEnablehscl000001r_ena <= '0' ;
      outp_ena <= '0' ;
      
      cond1_sT := 
      and2(bc_unsigned_ne(ihscl0000063,   conv_std_logic_vector(1,  10)),  bc_unsigned_lt
                                                                    (ihscl0000063,   conv_std_logic_vector
                                                                    (63,  10))) 
      ;
      h1_cond1sT_synchscl000006f <= cond1_sT ;
      tmp := 
      arrayTrim(sumsqshscl0000066,  conv_std_logic_vector(conv_std_logic_vector
                                                          (bc_unsigned_sub
                                                           (ihscl0000063,   conv_std_logic_vector
                                                                    (1,  10))))) 
      ;
      qssumsqs_sT := bc_unsigned_c_ext(tmp,  48) ;
      h1_qssumsqssT_synchscl000006g <= qssumsqs_sT ;
      tmp1 := 
      arrayTrim(sumshscl0000065,  conv_std_logic_vector(conv_std_logic_vector
                                                        (bc_unsigned_sub
                                                         (ihscl0000063,   conv_std_logic_vector
                                                                    (1,  10))))) 
      ;
      tmp2 := 
      arrayTrim(sumshscl0000065,  conv_std_logic_vector(conv_std_logic_vector
                                                        (bc_unsigned_sub
                                                         (ihscl0000063,   conv_std_logic_vector
                                                                    (1,  10))))) 
      ;
      qssums_sT := 
      conv_std_logic_vector(conv_std_logic_vector(bc_signed_emul(tmp1,  tmp2))) 
      ;
      h1_qssumssT_synchscl000006h <= qssums_sT ;
      tmp3 := 
      generic_std_logic_vector_trim(conv_std_logic_vector(shrConst(bc_unsigned_emul
                                                                   (qssumsqs_sT,  bc_unsigned_c_ext
                                                                    (arrayTrim
                                                                    (icoefmulthscl0000064,  ihscl0000063),  48)),  12)),  0,  63) 
      ;
      tmp4 := 
      bc_unsigned_c_ext(bc_unsigned_emul(arrayTrim(icoefmulthscl0000064,  ihscl0000063),  arrayTrim
                                                                    (icoefmulthscl0000064,  ihscl0000063)),  48) 
      ;
      tmp5 := 
       conv_std_logic_vector(generic_std_logic_vector_trim(conv_std_logic_vector
                                                           (shrConst(bc_unsigned_emul
                                                                    (qssums_sT,  tmp4),  24)),  0,  63)) 
      ;
      varL_sT := bc_unsigned_sub( conv_std_logic_vector(tmp3),  tmp5) ;
      h1_varLsT_synchscl000006i <= varL_sT ;
      
      cond_sT := equal(ihscl0000063,   conv_std_logic_vector(62,  10)) ;
      h1_condsT_synchscl000006j <= cond_sT ;
      
      null;
      
      outp_data <= 
      (p3 => endofoutphscl0000036,  p2 => varL_sT,  p1 => bc_unsigned_c_ext
                                                          (qssums_sT,  64),  p0 => bc_unsigned_c_ext
                                                                    (qssumsqs_sT,  64)) 
      ;
      
      null;
      
      null;
      
      h1sTTE_finish3hscl000001b_data <= 
      (p0 => h1sTTE_finish2hscl0000019_data.p0) ;
      
      null;
      h1sTET_cond_synchscl000006n_data_dummy := 
      zero(h1sTET_cond_synchscl000006n_data_dummy) ;
      h1sTET_cond_synchscl000006n <= h1sTET_cond_synchscl000006n_data_dummy ;
      h1sTE_cond_synchscl000006m_data_dummy := 
      zero(h1sTE_cond_synchscl000006m_data_dummy) ;
      h1sTE_cond_synchscl000006m <= h1sTE_cond_synchscl000006m_data_dummy ;
      h1sT_cond_synchscl000006k_data_dummy := 
      zero(h1sT_cond_synchscl000006k_data_dummy) ;
      h1sT_cond_synchscl000006k <= h1sT_cond_synchscl000006k_data_dummy ;
      h1s_cond_synchscl000006e_data_dummy := 
      zero(h1s_cond_synchscl000006e_data_dummy) ;
      h1s_cond_synchscl000006e <= h1s_cond_synchscl000006e_data_dummy ;
      h1sT_cond_sync1hscl000006l_data_dummy := 
      zero(h1sT_cond_sync1hscl000006l_data_dummy) ;
      h1sT_cond_sync1hscl000006l <= h1sT_cond_sync1hscl000006l_data_dummy ;
      
      s_condExpr := and2(not2((0 => '0')),  (0 => '1')) ;
      s_cond := (s_condExpr(0)) and h1sTTE_finish2hscl0000019_ena ;
      h1s_cond_synchscl000006e <= (0 => s_cond) ;
      if (s_cond='1') then
        h1_thenEnablehscl000001l_ena <= '1' ;
        null;
        h1_then_enablehscl000001m_ena <= '1' ;
        null;
        
        sT_condExpr5 := h1_then_leftHappenedhscl000003f ;
        sT_cond5 := (sT_condExpr5(0)) ;
        h1sT_cond_sync1hscl000006l <= (0 => sT_cond5) ;
        if (sT_cond5='1') then
          null;
        else
          
          sTE_condExpr := and2(not2((0 => '0')),  cond1_sT) ;
          sTE_cond := (sTE_condExpr(0)) ;
          h1sTE_cond_synchscl000006m <= (0 => sTE_cond) ;
          if (sTE_cond='1') then
            h1_then_l_thenEnablehscl000001o_ena <= '1' ;
            null;
            
            sTET_condExpr := and2(not2((0 => '0')),  cond_sT) ;
            sTET_cond := (sTET_condExpr(0)) ;
            h1sTET_cond_synchscl000006n <= (0 => sTET_cond) ;
            if (sTET_cond='1') then
              h1_then_l_then_p2_thenEnablehscl000001r_ena <= '1' ;
              null;
            else
              null;
            end if;
            outp_ena <= '1' ;
            null;
          else
            null;
          end if;
        end if;
        
        sT_condExpr := (0 => h1_then_rightEnablehscl000001s_ena) ;
        sT_cond := (sT_condExpr(0)) ;
        h1sT_cond_synchscl000006k <= (0 => sT_cond) ;
        if (sT_cond='1') then
          h1sTTE_finish3hscl000001b_ena <= '1' ;
          null;
        else
          null;
        end if;
      else
        null;
      end if;
      null;
    end process;
    process (h1sTTE_finish4hscl000001d_ena, h1sTTE_finish4hscl000001d_data, h1sTT_finishhscl000001t_ena, h1sTT_finishhscl000001t_data) 
    is
    variable s_condExpr : std_logic_vector (0 downto 0) ;
    variable s_cond : std_logic ;
    variable sE_condExpr : std_logic_vector (0 downto 0) ;
    variable sE_cond : std_logic ;
    variable h2sE_cond_synchscl000006p_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h2s_cond_synchscl000006o_data_dummy : 
    std_logic_vector (0 downto 0) ;
    begin
      h2_thenEnablehscl0000026_ena <= '0' ;
      h1sTT_finish4hscl000001u_ena <= '0' ;
      h2_else_thenEnablehscl0000025_ena <= '0' ;
      
      
      null;
      
      null;
      
      h1sTT_finish4hscl000001u_data <= 
      (p0 => h1sTT_finishhscl000001t_data.p0) ;
      h2s_cond_synchscl000006o_data_dummy := 
      zero(h2s_cond_synchscl000006o_data_dummy) ;
      h2s_cond_synchscl000006o <= h2s_cond_synchscl000006o_data_dummy ;
      h2sE_cond_synchscl000006p_data_dummy := 
      zero(h2sE_cond_synchscl000006p_data_dummy) ;
      h2sE_cond_synchscl000006p <= h2sE_cond_synchscl000006p_data_dummy ;
      
      s_condExpr := and2(not2((0 => '0')),  (0 => '1')) ;
      s_cond := (s_condExpr(0)) and h1sTT_finishhscl000001t_ena ;
      h2s_cond_synchscl000006o <= (0 => s_cond) ;
      if (s_cond='1') then
        h2_thenEnablehscl0000026_ena <= '1' ;
        null;
        h1sTT_finish4hscl000001u_ena <= '1' ;
        null;
      else
        
        sE_condExpr := and2(not2((0 => '0')),  (0 => '1')) ;
        sE_cond := (sE_condExpr(0)) and h1sTTE_finish4hscl000001d_ena ;
        h2sE_cond_synchscl000006p <= (0 => sE_cond) ;
        if (sE_cond='1') then
          h2_else_thenEnablehscl0000025_ena <= '1' ;
          null;
          h1sTT_finish4hscl000001u_ena <= '1' ;
          
          h1sTT_finish4hscl000001u_data <= 
          (p0 => h1sTTE_finish4hscl000001d_data.p0) ;
        else
          null;
        end if;
      end if;
      null;
    end process;
    process (h1sT_finishhscl000001x_ena, h1sTT_finish4hscl000001u_ena, h1sT_finishhscl000001x_data, h1sTT_finish4hscl000001u_data) 
    is
    variable s_condExpr : std_logic_vector (0 downto 0) ;
    variable s_cond : std_logic ;
    variable sE_condExpr : std_logic_vector (0 downto 0) ;
    variable sE_cond : std_logic ;
    variable h3s_cond_synchscl000006q_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h3sE_cond_synchscl000006r_data_dummy : 
    std_logic_vector (0 downto 0) ;
    begin
      h3_else_thenEnablehscl0000029_ena <= '0' ;
      h3_thenEnablehscl000002a_ena <= '0' ;
      h1sT_finish4hscl000001y_ena <= '0' ;
      
      
      null;
      
      h1sT_finish4hscl000001y_data <= 
      (p0 => h1sTT_finish4hscl000001u_data.p0) ;
      
      null;
      h3sE_cond_synchscl000006r_data_dummy := 
      zero(h3sE_cond_synchscl000006r_data_dummy) ;
      h3sE_cond_synchscl000006r <= h3sE_cond_synchscl000006r_data_dummy ;
      h3s_cond_synchscl000006q_data_dummy := 
      zero(h3s_cond_synchscl000006q_data_dummy) ;
      h3s_cond_synchscl000006q <= h3s_cond_synchscl000006q_data_dummy ;
      
      s_condExpr := and2(not2((0 => '0')),  (0 => '1')) ;
      s_cond := (s_condExpr(0)) and h1sTT_finish4hscl000001u_ena ;
      h3s_cond_synchscl000006q <= (0 => s_cond) ;
      if (s_cond='1') then
        h3_thenEnablehscl000002a_ena <= '1' ;
        null;
        h1sT_finish4hscl000001y_ena <= '1' ;
        null;
      else
        
        sE_condExpr := and2(not2((0 => '0')),  (0 => '1')) ;
        sE_cond := (sE_condExpr(0)) and h1sT_finishhscl000001x_ena ;
        h3sE_cond_synchscl000006r <= (0 => sE_cond) ;
        if (sE_cond='1') then
          h3_else_thenEnablehscl0000029_ena <= '1' ;
          null;
          h1sT_finish4hscl000001y_ena <= '1' ;
          
          h1sT_finish4hscl000001y_data <= 
          (p0 => h1sT_finishhscl000001x_data.p0) ;
        else
          null;
        end if;
      end if;
      null;
    end process;
    process (h1sT_finish4hscl000001y_data, h1sT_finish4hscl000001y_ena) is
    variable s_condExpr : std_logic_vector (0 downto 0) ;
    variable s_cond : std_logic ;
    variable h4s_cond_synchscl000006s_data_dummy : 
    std_logic_vector (0 downto 0) ;
    begin
      h4_thenEnablehscl000002c_ena <= '0' ;
      h1s_finish4hscl0000021_ena <= '0' ;
      
      
      null;
      
      null;
      h4s_cond_synchscl000006s_data_dummy := 
      zero(h4s_cond_synchscl000006s_data_dummy) ;
      h4s_cond_synchscl000006s <= h4s_cond_synchscl000006s_data_dummy ;
      
      s_condExpr := and2(not2((0 => '0')),  (0 => '1')) ;
      s_cond := (s_condExpr(0)) and h1sT_finish4hscl000001y_ena ;
      h4s_cond_synchscl000006s <= (0 => s_cond) ;
      if (s_cond='1') then
        h4_thenEnablehscl000002c_ena <= '1' ;
        null;
        h1s_finish4hscl0000021_ena <= '1' ;
        null;
      else
        null;
      end if;
      null;
    end process;
    process (inp_ena, sumshscl0000065, sumsqshscl0000066, h5_then_then_then_rightEnablehscl000002q_ena, reset_ena, h5_then_then_elseTransactionhscl000003n, h5_then_then_else_leftHappenedhscl000003s, inp_data, h5_then_then_then_leftHappenedhscl000003w, ihscl0000063, h5_then_then_else_rightEnablehscl000002m_ena) 
    is
    variable s_condExpr : std_logic_vector (0 downto 0) ;
    variable s_cond : std_logic ;
    variable sT_condExpr : std_logic_vector (0 downto 0) ;
    variable sT_cond : std_logic ;
    variable sTT_condExpr : std_logic_vector (0 downto 0) ;
    variable sTT_cond : std_logic ;
    variable sTTT_condExpr : std_logic_vector (0 downto 0) ;
    variable sTTT_cond : std_logic ;
    variable sTTT_condExpr1 : std_logic_vector (0 downto 0) ;
    variable sTTT_cond1 : std_logic ;
    variable cond_sTTE : std_logic_vector (0 downto 0) ;
    variable sTTE_condExpr : std_logic_vector (0 downto 0) ;
    variable sTTE_cond : std_logic ;
    variable sTTE_condExpr1 : std_logic_vector (0 downto 0) ;
    variable sTTE_cond1 : std_logic ;
    variable sTTEE_condExpr : std_logic_vector (0 downto 0) ;
    variable sTTEE_cond : std_logic ;
    variable h5sTTE_cond_sync1hscl0000070_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h5sTTT_cond_synchscl000006w_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h5sTTEE_cond_synchscl0000071_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h5sTTE_cond_synchscl000006z_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h5sTT_cond_synchscl000006v_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h5s_cond_synchscl000006t_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h5sT_cond_synchscl000006u_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h5sTTT_cond_sync1hscl000006x_data_dummy : 
    std_logic_vector (0 downto 0) ;
    begin
      h5_then_thenEnablehscl000002g_ena <= '0' ;
      h1sT_finishhscl000001x_ena <= '0' ;
      h5_thenEnablehscl000002e_ena <= '0' ;
      h1sTTE_finishhscl0000013_ena <= '0' ;
      h5_then_then_elseEnablehscl000002h_ena <= '0' ;
      h5_then_then_else_l_p0_thenEnablehscl000002l_ena <= '0' ;
      h5_then_then_then_enablehscl000002o_ena <= '0' ;
      h1sTT_finishhscl000001t_ena <= '0' ;
      h5_then_then_thenEnablehscl000002n_ena <= '0' ;
      h5_then_then_else_enablehscl000002i_ena <= '0' ;
      
      cond_sTTE := equal(ihscl0000063,   conv_std_logic_vector(63,  10)) ;
      h5_condsTTE_synchscl000006y <= cond_sTTE ;
      
      null;
      
      null;
      
      null;
      
      h1sT_finishhscl000001x_data <= (p0 => inp_data.p0) ;
      
      null;
      
      null;
      
      h1sTTE_finishhscl0000013_data <= (p0 => inp_data.p0) ;
      
      null;
      
      h1sTT_finishhscl000001t_data <= (p0 => inp_data.p0) ;
      
      null;
      h5sTTT_cond_sync1hscl000006x_data_dummy := 
      zero(h5sTTT_cond_sync1hscl000006x_data_dummy) ;
      h5sTTT_cond_sync1hscl000006x <= 
      h5sTTT_cond_sync1hscl000006x_data_dummy ;
      h5sT_cond_synchscl000006u_data_dummy := 
      zero(h5sT_cond_synchscl000006u_data_dummy) ;
      h5sT_cond_synchscl000006u <= h5sT_cond_synchscl000006u_data_dummy ;
      h5s_cond_synchscl000006t_data_dummy := 
      zero(h5s_cond_synchscl000006t_data_dummy) ;
      h5s_cond_synchscl000006t <= h5s_cond_synchscl000006t_data_dummy ;
      h5sTT_cond_synchscl000006v_data_dummy := 
      zero(h5sTT_cond_synchscl000006v_data_dummy) ;
      h5sTT_cond_synchscl000006v <= h5sTT_cond_synchscl000006v_data_dummy ;
      h5sTTE_cond_synchscl000006z_data_dummy := 
      zero(h5sTTE_cond_synchscl000006z_data_dummy) ;
      h5sTTE_cond_synchscl000006z <= h5sTTE_cond_synchscl000006z_data_dummy ;
      h5sTTEE_cond_synchscl0000071_data_dummy := 
      zero(h5sTTEE_cond_synchscl0000071_data_dummy) ;
      h5sTTEE_cond_synchscl0000071 <= 
      h5sTTEE_cond_synchscl0000071_data_dummy ;
      h5sTTT_cond_synchscl000006w_data_dummy := 
      zero(h5sTTT_cond_synchscl000006w_data_dummy) ;
      h5sTTT_cond_synchscl000006w <= h5sTTT_cond_synchscl000006w_data_dummy ;
      h5sTTE_cond_sync1hscl0000070_data_dummy := 
      zero(h5sTTE_cond_sync1hscl0000070_data_dummy) ;
      h5sTTE_cond_sync1hscl0000070 <= 
      h5sTTE_cond_sync1hscl0000070_data_dummy ;
      
      s_condExpr := 
      and2(not2((0 => '0')),  and2(not2((0 => reset_ena)),  (0 => '1'))) ;
      s_cond := (s_condExpr(0)) and inp_ena ;
      h5s_cond_synchscl000006t <= (0 => s_cond) ;
      if (s_cond='1') then
        h5_thenEnablehscl000002e_ena <= '1' ;
        null;
        
        sT_condExpr := 
        and2(not2((0 => '0')),  bc_unsigned_lt(ihscl0000063,   conv_std_logic_vector
                                                              (64,  10))) ;
        sT_cond := (sT_condExpr(0)) ;
        h5sT_cond_synchscl000006u <= (0 => sT_cond) ;
        if (sT_cond='1') then
          h5_then_thenEnablehscl000002g_ena <= '1' ;
          null;
          
          sTT_condExpr := 
          and2(not2(h5_then_then_elseTransactionhscl000003n),  equal(ihscl0000063,   conv_std_logic_vector
                                                                    (0,  10))) 
          ;
          sTT_cond := (sTT_condExpr(0)) ;
          h5sTT_cond_synchscl000006v <= (0 => sTT_cond) ;
          if (sTT_cond='1') then
            h5_then_then_thenEnablehscl000002n_ena <= '1' ;
            null;
            h5_then_then_then_enablehscl000002o_ena <= '1' ;
            null;
            
            sTTT_condExpr1 := h5_then_then_then_leftHappenedhscl000003w ;
            sTTT_cond1 := (sTTT_condExpr1(0)) ;
            h5sTTT_cond_sync1hscl000006x <= (0 => sTTT_cond1) ;
            if (sTTT_cond1='1') then
              null;
            else
              null;
            end if;
            
            sTTT_condExpr := 
            (0 => h5_then_then_then_rightEnablehscl000002q_ena) ;
            sTTT_cond := (sTTT_condExpr(0)) ;
            h5sTTT_cond_synchscl000006w <= (0 => sTTT_cond) ;
            if (sTTT_cond='1') then
              h1sTT_finishhscl000001t_ena <= '1' ;
              null;
            else
              null;
            end if;
          else
            h5_then_then_elseEnablehscl000002h_ena <= '1' ;
            null;
            h5_then_then_else_enablehscl000002i_ena <= '1' ;
            null;
            
            sTTE_condExpr1 := h5_then_then_else_leftHappenedhscl000003s ;
            sTTE_cond1 := (sTTE_condExpr1(0)) ;
            h5sTTE_cond_sync1hscl0000070 <= (0 => sTTE_cond1) ;
            if (sTTE_cond1='1') then
              null;
            else
              
              sTTEE_condExpr := and2(not2((0 => '0')),  cond_sTTE) ;
              sTTEE_cond := (sTTEE_condExpr(0)) ;
              h5sTTEE_cond_synchscl0000071 <= (0 => sTTEE_cond) ;
              if (sTTEE_cond='1') then
                h5_then_then_else_l_p0_thenEnablehscl000002l_ena <= '1' ;
                null;
              else
                null;
              end if;
            end if;
            
            sTTE_condExpr := 
            (0 => h5_then_then_else_rightEnablehscl000002m_ena) ;
            sTTE_cond := (sTTE_condExpr(0)) ;
            h5sTTE_cond_synchscl000006z <= (0 => sTTE_cond) ;
            if (sTTE_cond='1') then
              h1sTTE_finishhscl0000013_ena <= '1' ;
              null;
            else
              null;
            end if;
          end if;
        else
          h1sT_finishhscl000001x_ena <= '1' ;
          null;
        end if;
      else
        null;
      end if;
      null;
    end process;
    process (h1s_finish4hscl0000021_ena) is
    variable s_condExpr : std_logic_vector (0 downto 0) ;
    variable s_cond : std_logic ;
    variable h6s_cond_synchscl0000072_data_dummy : 
    std_logic_vector (0 downto 0) ;
    begin
      h6_thenEnablehscl000002s_ena <= '0' ;
      
      
      null;
      h6s_cond_synchscl0000072_data_dummy := 
      zero(h6s_cond_synchscl0000072_data_dummy) ;
      h6s_cond_synchscl0000072 <= h6s_cond_synchscl0000072_data_dummy ;
      
      s_condExpr := and2(not2((0 => '0')),  (0 => '1')) ;
      s_cond := (s_condExpr(0)) and h1s_finish4hscl0000021_ena ;
      h6s_cond_synchscl0000072 <= (0 => s_cond) ;
      if (s_cond='1') then
        h6_thenEnablehscl000002s_ena <= '1' ;
        null;
      else
        null;
      end if;
      null;
    end process;
    process (sumshscl0000065, varLefthscl0000067, sumsqshscl0000066, defihscl0000035, reset_ena, varRighthscl000006a, icoefmulthscl0000064, endofoutp1hscl0000037, ihscl0000063) 
    is
    variable s_condExpr : std_logic_vector (0 downto 0) ;
    variable s_cond : std_logic ;
    variable sT_condExpr : std_logic_vector (0 downto 0) ;
    variable sT_cond : std_logic ;
    variable subsumsqs_sTT :  std_logic_vector (48-1 downto 0) ;
    variable tmp :  std_logic_vector (32-1 downto 0) ;
    variable qssubsums_sTT :  std_logic_vector (48-1 downto 0) ;
    variable tmp1 :  std_logic_vector (24-1 downto 0) ;
    variable tmp2 :  std_logic_vector (24-1 downto 0) ;
    variable tmp3 :  std_logic_vector (48-1 downto 0) ;
    variable varR_sTT :  std_logic_vector (64-1 downto 0) ;
    variable tmp4 :  std_logic_vector (10-1 downto 0) ;
    variable tmp5 :  std_logic_vector (48-1 downto 0) ;
    variable tmp6 :  std_logic_vector (64-1 downto 0) ;
    variable tmp7 :  std_logic_vector (10-1 downto 0) ;
    variable tmp8 :  std_logic_vector (10-1 downto 0) ;
    variable tmp9 :  std_logic_vector (26-1 downto 0) ;
    variable tmp10 :  std_logic_vector (64-1 downto 0) ;
    variable tmp11 :  std_logic_vector (10-1 downto 0) ;
    variable tmp12 :  std_logic_vector (10-1 downto 0) ;
    variable sTT_condExpr : std_logic_vector (0 downto 0) ;
    variable sTT_cond : std_logic ;
    variable tmp13 : std_logic_vector (0 downto 0) ;
    variable sT_condExpr13 : std_logic_vector (0 downto 0) ;
    variable sT_cond13 : std_logic ;
    variable h7sTT_cond_synchscl0000078_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h7s_cond_synchscl0000073_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h7sT_cond_synchscl0000074_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h7sT_cond_sync1hscl0000079_data_dummy : 
    std_logic_vector (0 downto 0) ;
    begin
      outp1_ena <= '0' ;
      h7_then_p1_thenEnablehscl0000033_ena <= '0' ;
      h7_thenEnablehscl000002u_ena <= '0' ;
      outpVars_ena <= '0' ;
      h7_then_p0_then_p2_p2_thenEnablehscl0000031_ena <= '0' ;
      h7_then_p0_thenEnablehscl000002x_ena <= '0' ;
      tmp := 
      arrayTrim(sumsqshscl0000066,  conv_std_logic_vector(conv_std_logic_vector
                                                          (bc_unsigned_sub
                                                           (ihscl0000063,   conv_std_logic_vector
                                                                    (64,  10))))) 
      ;
      subsumsqs_sTT := 
      bc_unsigned_c_ext(bc_unsigned_sub(arrayTrim(sumsqshscl0000066,   conv_std_logic_vector
                                                                    (63,  10)),  tmp),  48) 
      ;
      h7_subsumsqssTT_synchscl0000075 <= subsumsqs_sTT ;
      tmp1 := 
      arrayTrim(sumshscl0000065,  conv_std_logic_vector(conv_std_logic_vector
                                                        (bc_unsigned_sub
                                                         (ihscl0000063,   conv_std_logic_vector
                                                                    (64,  10))))) 
      ;
      tmp2 := 
      arrayTrim(sumshscl0000065,  conv_std_logic_vector(conv_std_logic_vector
                                                        (bc_unsigned_sub
                                                         (ihscl0000063,   conv_std_logic_vector
                                                                    (64,  10))))) 
      ;
      tmp3 := 
      bc_signed_emul(bc_signed_sub(arrayTrim(sumshscl0000065,   conv_std_logic_vector
                                                               (63,  10)),  tmp1),  bc_signed_sub
                                                                    (arrayTrim
                                                                    (sumshscl0000065,   conv_std_logic_vector
                                                                    (63,  10)),  tmp2)) 
      ;
      qssubsums_sTT := conv_std_logic_vector(conv_std_logic_vector(tmp3)) ;
      h7_qssubsumssTT_synchscl0000076 <= qssubsums_sTT ;
      tmp4 := 
      bc_unsigned_sub( conv_std_logic_vector(64,  10),  bc_unsigned_sub
                                                        (bc_unsigned_add
                                                         (ihscl0000063,   conv_std_logic_vector
                                                                    (1,  10)),   conv_std_logic_vector
                                                                    (64,  10))) 
      ;
      tmp5 := 
      bc_unsigned_c_ext(arrayTrim(icoefmulthscl0000064,  conv_std_logic_vector
                                                         (conv_std_logic_vector
                                                          (tmp4))),  48) ;
      tmp6 := 
       conv_std_logic_vector(generic_std_logic_vector_trim(conv_std_logic_vector
                                                           (shrConst(bc_unsigned_emul
                                                                    (subsumsqs_sTT,  tmp5),  12)),  0,  63)) 
      ;
      tmp7 := 
      bc_unsigned_sub( conv_std_logic_vector(64,  10),  bc_unsigned_sub
                                                        (bc_unsigned_add
                                                         (ihscl0000063,   conv_std_logic_vector
                                                                    (1,  10)),   conv_std_logic_vector
                                                                    (64,  10))) 
      ;
      tmp8 := 
      bc_unsigned_sub( conv_std_logic_vector(64,  10),  bc_unsigned_sub
                                                        (bc_unsigned_add
                                                         (ihscl0000063,   conv_std_logic_vector
                                                                    (1,  10)),   conv_std_logic_vector
                                                                    (64,  10))) 
      ;
      tmp9 := 
      bc_unsigned_emul(arrayTrim(icoefmulthscl0000064,  conv_std_logic_vector
                                                        (conv_std_logic_vector
                                                         (tmp7))),  arrayTrim
                                                                    (icoefmulthscl0000064,  conv_std_logic_vector
                                                                    (conv_std_logic_vector
                                                                    (tmp8)))) 
      ;
      tmp10 := 
      generic_std_logic_vector_trim(conv_std_logic_vector(shrConst(bc_unsigned_emul
                                                                   (qssubsums_sTT,  bc_unsigned_c_ext
                                                                    (tmp9,  48)),  24)),  0,  63) 
      ;
      varR_sTT := bc_unsigned_sub(tmp6,   conv_std_logic_vector(tmp10)) ;
      h7_varRsTT_synchscl0000077 <= varR_sTT ;
      
      null;
      tmp11 := 
      bc_unsigned_sub(bc_unsigned_sub(ihscl0000063,   conv_std_logic_vector
                                                     (64,  10)),   conv_std_logic_vector
                                                                  (1,  10)) ;
      tmp12 := 
      bc_unsigned_sub(bc_unsigned_sub(ihscl0000063,   conv_std_logic_vector
                                                     (64,  10)),   conv_std_logic_vector
                                                                  (1,  10)) ;
      outpVars_data <= 
      (p2 => arrayTrim(varRighthscl000006a,  conv_std_logic_vector(conv_std_logic_vector
                                                                   (tmp11))),  p1 => arrayTrim
                                                                    (varLefthscl0000067,  conv_std_logic_vector
                                                                    (conv_std_logic_vector
                                                                    (tmp12))),  p0 => ihscl0000063) 
      ;
      
      outp1_data <= 
      (p3 => endofoutp1hscl0000037,  p2 => varR_sTT,  p1 => bc_unsigned_c_ext
                                                            (qssubsums_sTT,  64),  p0 => bc_unsigned_c_ext
                                                                    (subsumsqs_sTT,  64)) 
      ;
      
      null;
      
      null;
      
      null;
      h7sT_cond_sync1hscl0000079_data_dummy := 
      zero(h7sT_cond_sync1hscl0000079_data_dummy) ;
      h7sT_cond_sync1hscl0000079 <= h7sT_cond_sync1hscl0000079_data_dummy ;
      h7sT_cond_synchscl0000074_data_dummy := 
      zero(h7sT_cond_synchscl0000074_data_dummy) ;
      h7sT_cond_synchscl0000074 <= h7sT_cond_synchscl0000074_data_dummy ;
      h7s_cond_synchscl0000073_data_dummy := 
      zero(h7s_cond_synchscl0000073_data_dummy) ;
      h7s_cond_synchscl0000073 <= h7s_cond_synchscl0000073_data_dummy ;
      h7sTT_cond_synchscl0000078_data_dummy := 
      zero(h7sTT_cond_synchscl0000078_data_dummy) ;
      h7sTT_cond_synchscl0000078 <= h7sTT_cond_synchscl0000078_data_dummy ;
      
      s_condExpr := 
      and2(not2((0 => '0')),  and2(not2((0 => reset_ena)),  (0 => '1'))) ;
      s_cond := (s_condExpr(0)) ;
      h7s_cond_synchscl0000073 <= (0 => s_cond) ;
      if (s_cond='1') then
        h7_thenEnablehscl000002u_ena <= '1' ;
        null;
        
        sT_condExpr13 := and2(not2((0 => '0')),  defihscl0000035) ;
        sT_cond13 := (sT_condExpr13(0)) ;
        h7sT_cond_sync1hscl0000079 <= (0 => sT_cond13) ;
        if (sT_cond13='1') then
          h7_then_p1_thenEnablehscl0000033_ena <= '1' ;
          null;
        else
          null;
        end if;
        tmp13 := 
        and2(bc_unsigned_gt(ihscl0000063,   conv_std_logic_vector(64,  10)),  bc_unsigned_lt
                                                                    (ihscl0000063,   conv_std_logic_vector
                                                                    (126,  10))) 
        ;
        sT_condExpr := and2(not2((0 => '0')),  tmp13) ;
        sT_cond := (sT_condExpr(0)) ;
        h7sT_cond_synchscl0000074 <= (0 => sT_cond) ;
        if (sT_cond='1') then
          h7_then_p0_thenEnablehscl000002x_ena <= '1' ;
          null;
          
          sTT_condExpr := 
          and2(not2((0 => '0')),  equal(ihscl0000063,   conv_std_logic_vector
                                                       (125,  10))) ;
          sTT_cond := (sTT_condExpr(0)) ;
          h7sTT_cond_synchscl0000078 <= (0 => sTT_cond) ;
          if (sTT_cond='1') then
            h7_then_p0_then_p2_p2_thenEnablehscl0000031_ena <= '1' ;
            null;
          else
            null;
          end if;
          outp1_ena <= '1' ;
          null;
          outpVars_ena <= '1' ;
          null;
        else
          null;
        end if;
      else
        null;
      end if;
      null;
    end process;
    process (outp1_rdy_ena, h5_then_thenEnablehscl000002g_ena, h3_else_thenEnablehscl0000029_ena, h5_thenEnablehscl000002e_ena, h6_thenEnablehscl000002s_ena, h4_thenEnablehscl000002c_ena, h5_then_then_elseEnablehscl000002h_ena, h3_thenEnablehscl000002a_ena, reset_ena, h2_thenEnablehscl0000026_ena, h5_then_then_then_enablehscl000002o_ena, h5_then_then_elseTransactionhscl000003n, h1_then_enablehscl000001m_ena, h1_thenEnablehscl000001l_ena, Pipe_h1sTTE0BufFullhscl0000018_ena, h0_thenEnablehscl000001j_ena, h5_then_then_else_leftHappenedhscl000003s, h5_then_then_then_leftHappenedhscl000003w, h1_then_leftHappenedhscl000003f, h2_else_thenEnablehscl0000025_ena, h5_then_then_else_enablehscl000002i_ena, h5_then_then_thenEnablehscl000002n_ena, outpVars_rdy_ena, outp_rdy_ena) 
    is
    variable outpVars_rdy_s : std_logic_vector (0 downto 0) ;
    variable outp1_rdy_s : std_logic_vector (0 downto 0) ;
    variable outp_rdy_s : std_logic_vector (0 downto 0) ;
    variable h1s_finish4_rdy_s : std_logic_vector (0 downto 0) ;
    variable handlerForVarRCut_rdy_s : std_logic_vector (0 downto 0) ;
    variable h0_rdy_s : std_logic_vector (0 downto 0) ;
    variable tmp : std_logic_vector (0 downto 0) ;
    variable h4_then_rdy_s : std_logic_vector (0 downto 0) ;
    variable h1sT_finish4_rdy_s : std_logic_vector (0 downto 0) ;
    variable h4_rdy_s : std_logic_vector (0 downto 0) ;
    variable tmp1 : std_logic_vector (0 downto 0) ;
    variable h3_then_rdy_s : std_logic_vector (0 downto 0) ;
    variable h3_else_then_rdy_s : std_logic_vector (0 downto 0) ;
    variable h1sT_finish_rdy_s : std_logic_vector (0 downto 0) ;
    variable h3_else_rdy_s : std_logic_vector (0 downto 0) ;
    variable tmp2 : std_logic_vector (0 downto 0) ;
    variable h1sTT_finish4_rdy_s : std_logic_vector (0 downto 0) ;
    variable h3_rdy_s : std_logic_vector (0 downto 0) ;
    variable tmp3 : std_logic_vector (0 downto 0) ;
    variable h2_then_rdy_s : std_logic_vector (0 downto 0) ;
    variable h2_else_then_rdy_s : std_logic_vector (0 downto 0) ;
    variable h1sTTE_finish4_rdy_s : std_logic_vector (0 downto 0) ;
    variable h2_else_rdy_s : std_logic_vector (0 downto 0) ;
    variable tmp4 : std_logic_vector (0 downto 0) ;
    variable h1sTT_finish_rdy_s : std_logic_vector (0 downto 0) ;
    variable h2_rdy_s : std_logic_vector (0 downto 0) ;
    variable tmp5 : std_logic_vector (0 downto 0) ;
    variable h1_then_r_rdy_s : std_logic_vector (0 downto 0) ;
    variable h1_then_leftHappening_s : std_logic_vector (0 downto 0) ;
    variable h1_then_enableRight_s : std_logic_vector (0 downto 0) ;
    variable h1_then_rdy_s : std_logic_vector (0 downto 0) ;
    variable h1sTTE_finish2_rdy_s : std_logic_vector (0 downto 0) ;
    variable h1_rdy_s : std_logic_vector (0 downto 0) ;
    variable tmp6 : std_logic_vector (0 downto 0) ;
    variable h5_then_then_then_r_rdy_s : std_logic_vector (0 downto 0) ;
    variable h5_then_then_then_leftHappening_s : 
    std_logic_vector (0 downto 0) ;
    variable h5_then_then_then_enableRight_s : std_logic_vector (0 downto 0) 
    ;
    variable h5_then_then_then_rdy_s : std_logic_vector (0 downto 0) ;
    variable h5_then_then_else_r_rdy_s : std_logic_vector (0 downto 0) ;
    variable h5_then_then_else_leftHappening_s : 
    std_logic_vector (0 downto 0) ;
    variable h5_then_then_else_enableRight_s : std_logic_vector (0 downto 0) 
    ;
    variable h5_then_then_else_rdy_s : std_logic_vector (0 downto 0) ;
    variable h5_then_then_rdy_s : std_logic_vector (0 downto 0) ;
    variable tmp7 : std_logic_vector (0 downto 0) ;
    variable h5_then_else_rdy_s : std_logic_vector (0 downto 0) ;
    variable h5_then_rdy_s : std_logic_vector (0 downto 0) ;
    variable tmp8 : std_logic_vector (0 downto 0) ;
    variable inp_rdy_s : std_logic_vector (0 downto 0) ;
    variable h5_rdy_s : std_logic_vector (0 downto 0) ;
    variable tmp9 : std_logic_vector (0 downto 0) ;
    variable s_condExpr : std_logic_vector (0 downto 0) ;
    variable s_cond : std_logic ;
    variable s_condExpr9 : std_logic_vector (0 downto 0) ;
    variable s_cond9 : std_logic ;
    variable s_condExpr10 : std_logic_vector (0 downto 0) ;
    variable s_cond10 : std_logic ;
    variable s_condExpr11 : std_logic_vector (0 downto 0) ;
    variable s_cond11 : std_logic ;
    variable s_condExpr12 : std_logic_vector (0 downto 0) ;
    variable s_cond12 : std_logic ;
    variable s_condExpr13 : std_logic_vector (0 downto 0) ;
    variable s_cond13 : std_logic ;
    variable s_condExpr14 : std_logic_vector (0 downto 0) ;
    variable s_cond14 : std_logic ;
    variable s_condExpr15 : std_logic_vector (0 downto 0) ;
    variable s_cond15 : std_logic ;
    variable s_condExpr16 : std_logic_vector (0 downto 0) ;
    variable s_cond16 : std_logic ;
    variable s_condExpr17 : std_logic_vector (0 downto 0) ;
    variable s_cond17 : std_logic ;
    variable s_condExpr18 : std_logic_vector (0 downto 0) ;
    variable s_cond18 : std_logic ;
    variable s_condExpr19 : std_logic_vector (0 downto 0) ;
    variable s_cond19 : std_logic ;
    variable h8s_cond_sync2hscl000008g_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h8s_cond_sync7hscl000008l_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h8s_cond_sync1hscl000008f_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h8s_cond_sync6hscl000008k_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h8s_cond_sync9hscl000008n_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h8s_cond_sync10hscl000008o_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h8s_cond_synchscl000008e_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h8s_cond_sync5hscl000008j_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h8s_cond_sync3hscl000008h_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h8s_cond_sync11hscl000008p_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h8s_cond_sync4hscl000008i_data_dummy : 
    std_logic_vector (0 downto 0) ;
    variable h8s_cond_sync8hscl000008m_data_dummy : 
    std_logic_vector (0 downto 0) ;
    begin
      h1sTT_finish_rdyhscl000001w_ena <= '0' ;
      h1sTT_finish4_rdyhscl000001v_ena <= '0' ;
      handlerForVarRCut_rdyhscl000001e_ena <= '0' ;
      h5_then_then_then_rightEnablehscl000002q_ena <= '0' ;
      h1s_finish4_rdyhscl0000022_ena <= '0' ;
      h1sTTE_finish4_rdyhscl000001a_ena <= '0' ;
      inp_rdy_ena <= '0' ;
      h1_then_rightEnablehscl000001s_ena <= '0' ;
      h1sT_finish4_rdyhscl000001z_ena <= '0' ;
      h1sT_finish_rdyhscl0000020_ena <= '0' ;
      h1sTTE_finish2_rdyhscl0000017_ena <= '0' ;
      h5_then_then_else_rightEnablehscl000002m_ena <= '0' ;
      
      outpVars_rdy_s := (0 => outpVars_rdy_ena) ;
      h8_outpVars_rdys_synchscl000007a <= outpVars_rdy_s ;
      
      outp1_rdy_s := (0 => outp1_rdy_ena) ;
      h8_outp1_rdys_synchscl000007b <= outp1_rdy_s ;
      
      outp_rdy_s := (0 => outp_rdy_ena) ;
      h8_outp_rdys_synchscl000007c <= outp_rdy_s ;
      
      h1s_finish4_rdy_s := (0 => h6_thenEnablehscl000002s_ena) ;
      h8_h1s_finish4_rdys_synchscl000007d <= h1s_finish4_rdy_s ;
      
      handlerForVarRCut_rdy_s := (0 => h0_thenEnablehscl000001j_ena) ;
      h8_handlerForVarRCut_rdys_synchscl000007e <= handlerForVarRCut_rdy_s ;
      if conv_boolean((0 => h0_thenEnablehscl000001j_ena)) then
        tmp := (0 => '1') ;
      else
        tmp := (0 => '0') ;
      end if;
      h0_rdy_s := tmp ;
      h8_h0_rdys_synchscl000007f <= h0_rdy_s ;
      
      h4_then_rdy_s := h1s_finish4_rdy_s ;
      h8_h4_then_rdys_synchscl000007g <= h4_then_rdy_s ;
      
      h1sT_finish4_rdy_s := 
      and2(h4_then_rdy_s,  (0 => h4_thenEnablehscl000002c_ena)) ;
      h8_h1sT_finish4_rdys_synchscl000007h <= h1sT_finish4_rdy_s ;
      if conv_boolean((0 => h4_thenEnablehscl000002c_ena)) then
        tmp1 := h4_then_rdy_s ;
      else
        tmp1 := (0 => '1') ;
      end if;
      h4_rdy_s := tmp1 ;
      h8_h4_rdys_synchscl000007i <= h4_rdy_s ;
      
      h3_then_rdy_s := h1sT_finish4_rdy_s ;
      h8_h3_then_rdys_synchscl000007j <= h3_then_rdy_s ;
      
      h3_else_then_rdy_s := h1sT_finish4_rdy_s ;
      h8_h3_else_then_rdys_synchscl000007k <= h3_else_then_rdy_s ;
      
      h1sT_finish_rdy_s := 
      and2(h3_else_then_rdy_s,  (0 => h3_else_thenEnablehscl0000029_ena)) ;
      h8_h1sT_finish_rdys_synchscl000007l <= h1sT_finish_rdy_s ;
      if conv_boolean((0 => h3_else_thenEnablehscl0000029_ena)) then
        tmp2 := h3_else_then_rdy_s ;
      else
        tmp2 := (0 => '1') ;
      end if;
      h3_else_rdy_s := tmp2 ;
      h8_h3_else_rdys_synchscl000007m <= h3_else_rdy_s ;
      
      h1sTT_finish4_rdy_s := 
      and2(h3_then_rdy_s,  (0 => h3_thenEnablehscl000002a_ena)) ;
      h8_h1sTT_finish4_rdys_synchscl000007n <= h1sTT_finish4_rdy_s ;
      if conv_boolean((0 => h3_thenEnablehscl000002a_ena)) then
        tmp3 := h3_then_rdy_s ;
      else
        tmp3 := h3_else_rdy_s ;
      end if;
      h3_rdy_s := tmp3 ;
      h8_h3_rdys_synchscl000007o <= h3_rdy_s ;
      
      h2_then_rdy_s := h1sTT_finish4_rdy_s ;
      h8_h2_then_rdys_synchscl000007p <= h2_then_rdy_s ;
      
      h2_else_then_rdy_s := h1sTT_finish4_rdy_s ;
      h8_h2_else_then_rdys_synchscl000007q <= h2_else_then_rdy_s ;
      
      h1sTTE_finish4_rdy_s := 
      and2(h2_else_then_rdy_s,  (0 => h2_else_thenEnablehscl0000025_ena)) ;
      h8_h1sTTE_finish4_rdys_synchscl000007r <= h1sTTE_finish4_rdy_s ;
      if conv_boolean((0 => h2_else_thenEnablehscl0000025_ena)) then
        tmp4 := h2_else_then_rdy_s ;
      else
        tmp4 := (0 => '1') ;
      end if;
      h2_else_rdy_s := tmp4 ;
      h8_h2_else_rdys_synchscl000007s <= h2_else_rdy_s ;
      
      h1sTT_finish_rdy_s := 
      and2(h2_then_rdy_s,  (0 => h2_thenEnablehscl0000026_ena)) ;
      h8_h1sTT_finish_rdys_synchscl000007t <= h1sTT_finish_rdy_s ;
      if conv_boolean((0 => h2_thenEnablehscl0000026_ena)) then
        tmp5 := h2_then_rdy_s ;
      else
        tmp5 := h2_else_rdy_s ;
      end if;
      h2_rdy_s := tmp5 ;
      h8_h2_rdys_synchscl000007u <= h2_rdy_s ;
      
      h1_then_r_rdy_s := h1sTTE_finish4_rdy_s ;
      h8_h1_then_r_rdys_synchscl000007v <= h1_then_r_rdy_s ;
      
      h1_then_leftHappening_s := (0 => h1_then_enablehscl000001m_ena) ;
      h8_h1_then_leftHappenings_synchscl000007w <= h1_then_leftHappening_s ;
      
      h1_then_enableRight_s := 
      or2(h1_then_leftHappening_s,  h1_then_leftHappenedhscl000003f) ;
      h8_h1_then_enableRights_synchscl000007x <= h1_then_enableRight_s ;
      
      h1_then_rdy_s := and2(h1_then_enableRight_s,  h1_then_r_rdy_s) ;
      h8_h1_then_rdys_synchscl000007y <= h1_then_rdy_s ;
      
      h1sTTE_finish2_rdy_s := 
      and2(h1_then_rdy_s,  (0 => h1_thenEnablehscl000001l_ena)) ;
      h8_h1sTTE_finish2_rdys_synchscl000007z <= h1sTTE_finish2_rdy_s ;
      if conv_boolean((0 => h1_thenEnablehscl000001l_ena)) then
        tmp6 := h1_then_rdy_s ;
      else
        tmp6 := (0 => '1') ;
      end if;
      h1_rdy_s := tmp6 ;
      h8_h1_rdys_synchscl0000080 <= h1_rdy_s ;
      
      h5_then_then_then_r_rdy_s := h1sTT_finish_rdy_s ;
      h8_h5_then_then_then_r_rdys_synchscl0000081 <= 
      h5_then_then_then_r_rdy_s ;
      
      h5_then_then_then_leftHappening_s := 
      (0 => h5_then_then_then_enablehscl000002o_ena) ;
      h8_h5_then_then_then_leftHappenings_synchscl0000082 <= 
      h5_then_then_then_leftHappening_s ;
      
      h5_then_then_then_enableRight_s := 
      or2(h5_then_then_then_leftHappening_s,  h5_then_then_then_leftHappenedhscl000003w) 
      ;
      h8_h5_then_then_then_enableRights_synchscl0000083 <= 
      h5_then_then_then_enableRight_s ;
      
      h5_then_then_then_rdy_s := 
      and2(h5_then_then_then_enableRight_s,  h5_then_then_then_r_rdy_s) ;
      h8_h5_then_then_then_rdys_synchscl0000084 <= h5_then_then_then_rdy_s ;
      
      h5_then_then_else_r_rdy_s := 
      or2(h1sTTE_finish2_rdy_s,  not2((0 => Pipe_h1sTTE0BufFullhscl0000018_ena))) 
      ;
      h8_h5_then_then_else_r_rdys_synchscl0000085 <= 
      h5_then_then_else_r_rdy_s ;
      
      h5_then_then_else_leftHappening_s := 
      (0 => h5_then_then_else_enablehscl000002i_ena) ;
      h8_h5_then_then_else_leftHappenings_synchscl0000086 <= 
      h5_then_then_else_leftHappening_s ;
      
      h5_then_then_else_enableRight_s := 
      or2(h5_then_then_else_leftHappening_s,  h5_then_then_else_leftHappenedhscl000003s) 
      ;
      h8_h5_then_then_else_enableRights_synchscl0000087 <= 
      h5_then_then_else_enableRight_s ;
      
      h5_then_then_else_rdy_s := 
      and2(h5_then_then_else_enableRight_s,  h5_then_then_else_r_rdy_s) ;
      h8_h5_then_then_else_rdys_synchscl0000088 <= h5_then_then_else_rdy_s ;
      if conv_boolean((0 => h5_then_then_thenEnablehscl000002n_ena)) then
        tmp7 := h5_then_then_then_rdy_s ;
      else
        tmp7 := h5_then_then_else_rdy_s ;
      end if;
      h5_then_then_rdy_s := tmp7 ;
      h8_h5_then_then_rdys_synchscl0000089 <= h5_then_then_rdy_s ;
      
      h5_then_else_rdy_s := h1sT_finish_rdy_s ;
      h8_h5_then_else_rdys_synchscl000008a <= h5_then_else_rdy_s ;
      if conv_boolean((0 => h5_then_thenEnablehscl000002g_ena)) then
        tmp8 := h5_then_then_rdy_s ;
      else
        tmp8 := h5_then_else_rdy_s ;
      end if;
      h5_then_rdy_s := tmp8 ;
      h8_h5_then_rdys_synchscl000008b <= h5_then_rdy_s ;
      
      inp_rdy_s := and2(h5_then_rdy_s,  (0 => h5_thenEnablehscl000002e_ena)) 
      ;
      h8_inp_rdys_synchscl000008c <= inp_rdy_s ;
      if conv_boolean((0 => h5_thenEnablehscl000002e_ena)) then
        tmp9 := h5_then_rdy_s ;
      else
        tmp9 := (0 => '0') ;
      end if;
      h5_rdy_s := tmp9 ;
      h8_h5_rdys_synchscl000008d <= h5_rdy_s ;
      
      null;
      
      null;
      
      null;
      
      null;
      
      null;
      
      null;
      
      null;
      
      null;
      
      null;
      
      null;
      
      null;
      
      null;
      h8s_cond_sync8hscl000008m_data_dummy := 
      zero(h8s_cond_sync8hscl000008m_data_dummy) ;
      h8s_cond_sync8hscl000008m <= h8s_cond_sync8hscl000008m_data_dummy ;
      h8s_cond_sync4hscl000008i_data_dummy := 
      zero(h8s_cond_sync4hscl000008i_data_dummy) ;
      h8s_cond_sync4hscl000008i <= h8s_cond_sync4hscl000008i_data_dummy ;
      h8s_cond_sync11hscl000008p_data_dummy := 
      zero(h8s_cond_sync11hscl000008p_data_dummy) ;
      h8s_cond_sync11hscl000008p <= h8s_cond_sync11hscl000008p_data_dummy ;
      h8s_cond_sync3hscl000008h_data_dummy := 
      zero(h8s_cond_sync3hscl000008h_data_dummy) ;
      h8s_cond_sync3hscl000008h <= h8s_cond_sync3hscl000008h_data_dummy ;
      h8s_cond_sync5hscl000008j_data_dummy := 
      zero(h8s_cond_sync5hscl000008j_data_dummy) ;
      h8s_cond_sync5hscl000008j <= h8s_cond_sync5hscl000008j_data_dummy ;
      h8s_cond_synchscl000008e_data_dummy := 
      zero(h8s_cond_synchscl000008e_data_dummy) ;
      h8s_cond_synchscl000008e <= h8s_cond_synchscl000008e_data_dummy ;
      h8s_cond_sync10hscl000008o_data_dummy := 
      zero(h8s_cond_sync10hscl000008o_data_dummy) ;
      h8s_cond_sync10hscl000008o <= h8s_cond_sync10hscl000008o_data_dummy ;
      h8s_cond_sync9hscl000008n_data_dummy := 
      zero(h8s_cond_sync9hscl000008n_data_dummy) ;
      h8s_cond_sync9hscl000008n <= h8s_cond_sync9hscl000008n_data_dummy ;
      h8s_cond_sync6hscl000008k_data_dummy := 
      zero(h8s_cond_sync6hscl000008k_data_dummy) ;
      h8s_cond_sync6hscl000008k <= h8s_cond_sync6hscl000008k_data_dummy ;
      h8s_cond_sync1hscl000008f_data_dummy := 
      zero(h8s_cond_sync1hscl000008f_data_dummy) ;
      h8s_cond_sync1hscl000008f <= h8s_cond_sync1hscl000008f_data_dummy ;
      h8s_cond_sync7hscl000008l_data_dummy := 
      zero(h8s_cond_sync7hscl000008l_data_dummy) ;
      h8s_cond_sync7hscl000008l <= h8s_cond_sync7hscl000008l_data_dummy ;
      h8s_cond_sync2hscl000008g_data_dummy := 
      zero(h8s_cond_sync2hscl000008g_data_dummy) ;
      h8s_cond_sync2hscl000008g <= h8s_cond_sync2hscl000008g_data_dummy ;
      
      s_condExpr19 := (0 => h6_thenEnablehscl000002s_ena) ;
      s_cond19 := (s_condExpr19(0)) ;
      h8s_cond_sync11hscl000008p <= (0 => s_cond19) ;
      if (s_cond19='1') then
        h1s_finish4_rdyhscl0000022_ena <= '1' ;
        null;
      else
        null;
      end if;
      
      s_condExpr18 := (0 => h0_thenEnablehscl000001j_ena) ;
      s_cond18 := (s_condExpr18(0)) ;
      h8s_cond_sync10hscl000008o <= (0 => s_cond18) ;
      if (s_cond18='1') then
        handlerForVarRCut_rdyhscl000001e_ena <= '1' ;
        null;
      else
        null;
      end if;
      
      s_condExpr17 := 
      and2(h4_then_rdy_s,  (0 => h4_thenEnablehscl000002c_ena)) ;
      s_cond17 := (s_condExpr17(0)) ;
      h8s_cond_sync9hscl000008n <= (0 => s_cond17) ;
      if (s_cond17='1') then
        h1sT_finish4_rdyhscl000001z_ena <= '1' ;
        null;
      else
        null;
      end if;
      
      s_condExpr16 := 
      and2(h3_else_then_rdy_s,  (0 => h3_else_thenEnablehscl0000029_ena)) ;
      s_cond16 := (s_condExpr16(0)) ;
      h8s_cond_sync8hscl000008m <= (0 => s_cond16) ;
      if (s_cond16='1') then
        h1sT_finish_rdyhscl0000020_ena <= '1' ;
        null;
      else
        null;
      end if;
      
      s_condExpr15 := 
      and2(h3_then_rdy_s,  (0 => h3_thenEnablehscl000002a_ena)) ;
      s_cond15 := (s_condExpr15(0)) ;
      h8s_cond_sync7hscl000008l <= (0 => s_cond15) ;
      if (s_cond15='1') then
        h1sTT_finish4_rdyhscl000001v_ena <= '1' ;
        null;
      else
        null;
      end if;
      
      s_condExpr14 := 
      and2(h2_else_then_rdy_s,  (0 => h2_else_thenEnablehscl0000025_ena)) ;
      s_cond14 := (s_condExpr14(0)) ;
      h8s_cond_sync6hscl000008k <= (0 => s_cond14) ;
      if (s_cond14='1') then
        h1sTTE_finish4_rdyhscl000001a_ena <= '1' ;
        null;
      else
        null;
      end if;
      
      s_condExpr13 := 
      and2(h2_then_rdy_s,  (0 => h2_thenEnablehscl0000026_ena)) ;
      s_cond13 := (s_condExpr13(0)) ;
      h8s_cond_sync5hscl000008j <= (0 => s_cond13) ;
      if (s_cond13='1') then
        h1sTT_finish_rdyhscl000001w_ena <= '1' ;
        null;
      else
        null;
      end if;
      
      s_condExpr12 := h1_then_enableRight_s ;
      s_cond12 := (s_condExpr12(0)) ;
      h8s_cond_sync4hscl000008i <= (0 => s_cond12) ;
      if (s_cond12='1') then
        h1_then_rightEnablehscl000001s_ena <= '1' ;
        null;
      else
        null;
      end if;
      
      s_condExpr11 := 
      and2(h1_then_rdy_s,  (0 => h1_thenEnablehscl000001l_ena)) ;
      s_cond11 := (s_condExpr11(0)) ;
      h8s_cond_sync3hscl000008h <= (0 => s_cond11) ;
      if (s_cond11='1') then
        h1sTTE_finish2_rdyhscl0000017_ena <= '1' ;
        null;
      else
        null;
      end if;
      
      s_condExpr10 := h5_then_then_then_enableRight_s ;
      s_cond10 := (s_condExpr10(0)) ;
      h8s_cond_sync2hscl000008g <= (0 => s_cond10) ;
      if (s_cond10='1') then
        h5_then_then_then_rightEnablehscl000002q_ena <= '1' ;
        null;
      else
        null;
      end if;
      
      s_condExpr9 := h5_then_then_else_enableRight_s ;
      s_cond9 := (s_condExpr9(0)) ;
      h8s_cond_sync1hscl000008f <= (0 => s_cond9) ;
      if (s_cond9='1') then
        h5_then_then_else_rightEnablehscl000002m_ena <= '1' ;
        null;
      else
        null;
      end if;
      
      s_condExpr := 
      and2(h5_then_rdy_s,  (0 => h5_thenEnablehscl000002e_ena)) ;
      s_cond := (s_condExpr(0)) ;
      h8s_cond_synchscl000008e <= (0 => s_cond) ;
      if (s_cond='1') then
        inp_rdy_ena <= '1' ;
        null;
      else
        null;
      end if;
      null;
    end process;
    process  is
    
    begin
      Pipe_h1sTTE0BufFull_rdyhscl0000016_ena <= '0' ;
      
      
      null;
      
      Pipe_h1sTTE0BufFull_rdyhscl0000016_ena <= '1' ;
      null;
      wait until false;
    end process;
    handlerForVarhscl000001f_ena <= '0' ;
    h7_then_p1_then_enablehscl0000034_ena <= '0' ;
    h7_then_p1_elseEnablehscl0000032_ena <= '0' ;
    h7_then_p0_then_p2_p2_elseEnablehscl0000030_ena <= '0' ;
    h7_then_p0_then_p2_enablehscl000002z_ena <= '0' ;
    h7_then_p0_then_enablehscl000002y_ena <= '0' ;
    h7_then_p0_elseEnablehscl000002w_ena <= '0' ;
    h7_then_enablehscl000002v_ena <= '0' ;
    h7_elseEnablehscl000002t_ena <= '0' ;
    h6_elseEnablehscl000002r_ena <= '0' ;
    h5_then_then_then_l_enablehscl000002p_ena <= '0' ;
    h5_then_then_else_l_p0_elseEnablehscl000002k_ena <= '0' ;
    h5_then_then_else_l_enablehscl000002j_ena <= '0' ;
    h5_then_elseEnablehscl000002f_ena <= '0' ;
    h5_elseEnablehscl000002d_ena <= '0' ;
    h4_elseEnablehscl000002b_ena <= '0' ;
    h3_else_elseEnablehscl0000028_ena <= '0' ;
    h3_elseEnablehscl0000027_ena <= '0' ;
    h2_else_elseEnablehscl0000024_ena <= '0' ;
    h2_elseEnablehscl0000023_ena <= '0' ;
    h1_then_l_then_p2_elseEnablehscl000001q_ena <= '0' ;
    h1_then_l_then_enablehscl000001p_ena <= '0' ;
    h1_then_l_elseEnablehscl000001n_ena <= '0' ;
    h1_elseEnablehscl000001k_ena <= '0' ;
    h0_elseEnablehscl000001i_ena <= '0' ;
    
end architecture;