library ieee;
use ieee.std_logic_1164.all;
library work;
use work.runtime.all;
package arrayAsAliasTrimmers is
  
end package;
package body arrayAsAliasTrimmers is 

end arrayAsAliasTrimmers;